
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_M32_C4_N5 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_M32_C4_N5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n11, n12 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n11, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n11);
   U1 : INV_X1 port map( A => n12, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n11, B2 => Ci, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_15;

architecture SYN_STRUCTURAL of RCA_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_14;

architecture SYN_STRUCTURAL of RCA_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_13;

architecture SYN_STRUCTURAL of RCA_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_12;

architecture SYN_STRUCTURAL of RCA_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_11;

architecture SYN_STRUCTURAL of RCA_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_10;

architecture SYN_STRUCTURAL of RCA_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_9;

architecture SYN_STRUCTURAL of RCA_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_8;

architecture SYN_STRUCTURAL of RCA_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_7;

architecture SYN_STRUCTURAL of RCA_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_6;

architecture SYN_STRUCTURAL of RCA_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_5;

architecture SYN_STRUCTURAL of RCA_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_4;

architecture SYN_STRUCTURAL of RCA_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_3;

architecture SYN_STRUCTURAL of RCA_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_2;

architecture SYN_STRUCTURAL of RCA_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_1;

architecture SYN_STRUCTURAL of RCA_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSb_6 is

   port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : out 
         std_logic_vector (3 downto 0));

end CSb_6;

architecture SYN_STRUCTURAL of CSb_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, 
      out0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, n26, n27
      , n28, n29, n30, n_1000, n_1001 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => out0_3_port, 
                           S(2) => out0_2_port, S(1) => out0_1_port, S(0) => 
                           out0_0_port, Co => n_1000);
   RCA1 : RCA_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => out1_3_port, 
                           S(2) => out1_2_port, S(1) => out1_1_port, S(0) => 
                           out1_0_port, Co => n_1001);
   U3 : INV_X1 port map( A => n30, ZN => s(3));
   U4 : INV_X1 port map( A => n29, ZN => s(2));
   U5 : INV_X1 port map( A => n28, ZN => s(1));
   U6 : INV_X1 port map( A => n27, ZN => s(0));
   U7 : AOI22_X1 port map( A1 => out0_3_port, A2 => n26, B1 => out1_3_port, B2 
                           => ci, ZN => n30);
   U8 : AOI22_X1 port map( A1 => out0_0_port, A2 => n26, B1 => out1_0_port, B2 
                           => ci, ZN => n27);
   U9 : AOI22_X1 port map( A1 => out0_1_port, A2 => n26, B1 => out1_1_port, B2 
                           => ci, ZN => n28);
   U10 : AOI22_X1 port map( A1 => out0_2_port, A2 => n26, B1 => out1_2_port, B2
                           => ci, ZN => n29);
   U11 : INV_X1 port map( A => ci, ZN => n26);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSb_5 is

   port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : out 
         std_logic_vector (3 downto 0));

end CSb_5;

architecture SYN_STRUCTURAL of CSb_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, 
      out0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, n26, n27
      , n28, n29, n30, n_1002, n_1003 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => out0_3_port, 
                           S(2) => out0_2_port, S(1) => out0_1_port, S(0) => 
                           out0_0_port, Co => n_1002);
   RCA1 : RCA_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => out1_3_port, 
                           S(2) => out1_2_port, S(1) => out1_1_port, S(0) => 
                           out1_0_port, Co => n_1003);
   U3 : INV_X1 port map( A => ci, ZN => n26);
   U4 : INV_X1 port map( A => n28, ZN => s(1));
   U5 : AOI22_X1 port map( A1 => out0_1_port, A2 => n26, B1 => out1_1_port, B2 
                           => ci, ZN => n28);
   U6 : INV_X1 port map( A => n29, ZN => s(2));
   U7 : AOI22_X1 port map( A1 => out0_2_port, A2 => n26, B1 => out1_2_port, B2 
                           => ci, ZN => n29);
   U8 : INV_X1 port map( A => n30, ZN => s(3));
   U9 : AOI22_X1 port map( A1 => out0_3_port, A2 => n26, B1 => out1_3_port, B2 
                           => ci, ZN => n30);
   U10 : INV_X1 port map( A => n27, ZN => s(0));
   U11 : AOI22_X1 port map( A1 => out0_0_port, A2 => n26, B1 => out1_0_port, B2
                           => ci, ZN => n27);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSb_4 is

   port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : out 
         std_logic_vector (3 downto 0));

end CSb_4;

architecture SYN_STRUCTURAL of CSb_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, 
      out0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, n26, n27
      , n28, n29, n30, n_1004, n_1005 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => out0_3_port, 
                           S(2) => out0_2_port, S(1) => out0_1_port, S(0) => 
                           out0_0_port, Co => n_1004);
   RCA1 : RCA_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => out1_3_port, 
                           S(2) => out1_2_port, S(1) => out1_1_port, S(0) => 
                           out1_0_port, Co => n_1005);
   U3 : INV_X1 port map( A => n30, ZN => s(3));
   U4 : INV_X1 port map( A => n29, ZN => s(2));
   U5 : INV_X1 port map( A => n28, ZN => s(1));
   U6 : INV_X1 port map( A => n27, ZN => s(0));
   U7 : AOI22_X1 port map( A1 => out0_3_port, A2 => n26, B1 => out1_3_port, B2 
                           => ci, ZN => n30);
   U8 : AOI22_X1 port map( A1 => out0_2_port, A2 => n26, B1 => out1_2_port, B2 
                           => ci, ZN => n29);
   U9 : AOI22_X1 port map( A1 => out0_1_port, A2 => n26, B1 => out1_1_port, B2 
                           => ci, ZN => n28);
   U10 : AOI22_X1 port map( A1 => out0_0_port, A2 => n26, B1 => out1_0_port, B2
                           => ci, ZN => n27);
   U11 : INV_X1 port map( A => ci, ZN => n26);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSb_3 is

   port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : out 
         std_logic_vector (3 downto 0));

end CSb_3;

architecture SYN_STRUCTURAL of CSb_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component RCA_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, 
      out0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, n26, n27
      , n28, n29, n_1006, n_1007 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => out0_3_port, 
                           S(2) => out0_2_port, S(1) => out0_1_port, S(0) => 
                           out0_0_port, Co => n_1006);
   RCA1 : RCA_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => out1_3_port, 
                           S(2) => out1_2_port, S(1) => out1_1_port, S(0) => 
                           out1_0_port, Co => n_1007);
   U3 : MUX2_X1 port map( A => out0_1_port, B => out1_1_port, S => ci, Z => 
                           s(1));
   U4 : INV_X1 port map( A => n27, ZN => s(0));
   U5 : AOI22_X1 port map( A1 => out0_3_port, A2 => n26, B1 => out1_3_port, B2 
                           => ci, ZN => n29);
   U6 : AOI22_X1 port map( A1 => out0_2_port, A2 => n26, B1 => out1_2_port, B2 
                           => ci, ZN => n28);
   U7 : AOI22_X1 port map( A1 => out0_0_port, A2 => n26, B1 => out1_0_port, B2 
                           => ci, ZN => n27);
   U8 : INV_X1 port map( A => ci, ZN => n26);
   U9 : INV_X1 port map( A => n28, ZN => s(2));
   U10 : INV_X1 port map( A => n29, ZN => s(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSb_2 is

   port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : out 
         std_logic_vector (3 downto 0));

end CSb_2;

architecture SYN_STRUCTURAL of CSb_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, 
      out0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, n26, n27
      , n28, n29, n30, n_1008, n_1009 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => out0_3_port, 
                           S(2) => out0_2_port, S(1) => out0_1_port, S(0) => 
                           out0_0_port, Co => n_1008);
   RCA1 : RCA_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => out1_3_port, 
                           S(2) => out1_2_port, S(1) => out1_1_port, S(0) => 
                           out1_0_port, Co => n_1009);
   U3 : AOI22_X1 port map( A1 => out0_3_port, A2 => n26, B1 => out1_3_port, B2 
                           => ci, ZN => n30);
   U4 : AOI22_X1 port map( A1 => out0_2_port, A2 => n26, B1 => out1_2_port, B2 
                           => ci, ZN => n29);
   U5 : AOI22_X1 port map( A1 => out0_1_port, A2 => n26, B1 => out1_1_port, B2 
                           => ci, ZN => n28);
   U6 : AOI22_X1 port map( A1 => out0_0_port, A2 => n26, B1 => out1_0_port, B2 
                           => ci, ZN => n27);
   U7 : INV_X1 port map( A => ci, ZN => n26);
   U8 : INV_X1 port map( A => n29, ZN => s(2));
   U9 : INV_X1 port map( A => n28, ZN => s(1));
   U10 : INV_X1 port map( A => n27, ZN => s(0));
   U11 : INV_X1 port map( A => n30, ZN => s(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSb_1 is

   port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : out 
         std_logic_vector (3 downto 0));

end CSb_1;

architecture SYN_STRUCTURAL of CSb_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, 
      out0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, n26, n27
      , n28, n29, n30, n_1010, n_1011 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => out0_3_port, 
                           S(2) => out0_2_port, S(1) => out0_1_port, S(0) => 
                           out0_0_port, Co => n_1010);
   RCA1 : RCA_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => out1_3_port, 
                           S(2) => out1_2_port, S(1) => out1_1_port, S(0) => 
                           out1_0_port, Co => n_1011);
   U3 : AOI22_X1 port map( A1 => out0_3_port, A2 => n26, B1 => out1_3_port, B2 
                           => ci, ZN => n30);
   U4 : AOI22_X1 port map( A1 => out0_2_port, A2 => n26, B1 => out1_2_port, B2 
                           => ci, ZN => n29);
   U5 : AOI22_X1 port map( A1 => out0_1_port, A2 => n26, B1 => out1_1_port, B2 
                           => ci, ZN => n28);
   U6 : AOI22_X1 port map( A1 => out0_0_port, A2 => n26, B1 => out1_0_port, B2 
                           => ci, ZN => n27);
   U7 : INV_X1 port map( A => ci, ZN => n26);
   U8 : INV_X1 port map( A => n27, ZN => s(0));
   U9 : INV_X1 port map( A => n28, ZN => s(1));
   U10 : INV_X1 port map( A => n29, ZN => s(2));
   U11 : INV_X1 port map( A => n30, ZN => s(3));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_9 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_9;

architecture SYN_BEHAVIORAL of G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_8 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_8;

architecture SYN_BEHAVIORAL of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_7 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_7;

architecture SYN_BEHAVIORAL of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_6 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_6;

architecture SYN_BEHAVIORAL of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_5 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_5;

architecture SYN_BEHAVIORAL of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X2 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_4 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_4;

architecture SYN_BEHAVIORAL of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_3 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_3;

architecture SYN_BEHAVIORAL of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_2 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_2;

architecture SYN_BEHAVIORAL of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_1 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_1;

architecture SYN_BEHAVIORAL of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_30 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_30;

architecture SYN_BEHAVIORAL of PGnet_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_29 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_29;

architecture SYN_BEHAVIORAL of PGnet_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_28 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_28;

architecture SYN_BEHAVIORAL of PGnet_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_27 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_27;

architecture SYN_BEHAVIORAL of PGnet_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_26 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_26;

architecture SYN_BEHAVIORAL of PGnet_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_25 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_25;

architecture SYN_BEHAVIORAL of PGnet_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_24 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_24;

architecture SYN_BEHAVIORAL of PGnet_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_23 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_23;

architecture SYN_BEHAVIORAL of PGnet_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_22 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_22;

architecture SYN_BEHAVIORAL of PGnet_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_21 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_21;

architecture SYN_BEHAVIORAL of PGnet_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_20 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_20;

architecture SYN_BEHAVIORAL of PGnet_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_19 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_19;

architecture SYN_BEHAVIORAL of PGnet_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_18 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_18;

architecture SYN_BEHAVIORAL of PGnet_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_17 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_17;

architecture SYN_BEHAVIORAL of PGnet_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_16 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_16;

architecture SYN_BEHAVIORAL of PGnet_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_15 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_15;

architecture SYN_BEHAVIORAL of PGnet_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_14 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_14;

architecture SYN_BEHAVIORAL of PGnet_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_13 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_13;

architecture SYN_BEHAVIORAL of PGnet_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_12 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_12;

architecture SYN_BEHAVIORAL of PGnet_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_11 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_11;

architecture SYN_BEHAVIORAL of PGnet_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_10 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_10;

architecture SYN_BEHAVIORAL of PGnet_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_9 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_9;

architecture SYN_BEHAVIORAL of PGnet_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_8 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_8;

architecture SYN_BEHAVIORAL of PGnet_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_7 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_7;

architecture SYN_BEHAVIORAL of PGnet_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_6 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_6;

architecture SYN_BEHAVIORAL of PGnet_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_5 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_5;

architecture SYN_BEHAVIORAL of PGnet_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U3 : AND2_X1 port map( A1 => n1, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_4 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_4;

architecture SYN_BEHAVIORAL of PGnet_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_3 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_3;

architecture SYN_BEHAVIORAL of PGnet_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_2 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_2;

architecture SYN_BEHAVIORAL of PGnet_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_1 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_1;

architecture SYN_BEHAVIORAL of PGnet_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_8 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_8;

architecture SYN_behavioral of reg_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180, n181, n182,
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n215, Z => n177);
   U4 : BUF_X1 port map( A => n215, Z => n176);
   U5 : BUF_X1 port map( A => n215, Z => n178);
   U6 : BUF_X1 port map( A => n216, Z => n179);
   U7 : BUF_X1 port map( A => n216, Z => n180);
   U8 : BUF_X1 port map( A => n216, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n215);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U11 : INV_X1 port map( A => i(1), ZN => n213);
   U12 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U13 : INV_X1 port map( A => i(2), ZN => n212);
   U14 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U15 : INV_X1 port map( A => i(6), ZN => n208);
   U16 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U17 : INV_X1 port map( A => i(7), ZN => n207);
   U18 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U19 : INV_X1 port map( A => i(8), ZN => n206);
   U20 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U21 : INV_X1 port map( A => i(10), ZN => n204);
   U22 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U23 : INV_X1 port map( A => i(11), ZN => n203);
   U24 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U25 : INV_X1 port map( A => i(12), ZN => n202);
   U26 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U27 : INV_X1 port map( A => i(13), ZN => n201);
   U28 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U29 : INV_X1 port map( A => i(14), ZN => n200);
   U30 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n199, ZN 
                           => n84);
   U31 : INV_X1 port map( A => i(15), ZN => n199);
   U32 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n198, ZN 
                           => n83);
   U33 : INV_X1 port map( A => i(16), ZN => n198);
   U34 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n197, ZN 
                           => n82);
   U35 : INV_X1 port map( A => i(17), ZN => n197);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n196, ZN 
                           => n81);
   U37 : INV_X1 port map( A => i(18), ZN => n196);
   U38 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n195, ZN 
                           => n80);
   U39 : INV_X1 port map( A => i(19), ZN => n195);
   U40 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n194, ZN 
                           => n79);
   U41 : INV_X1 port map( A => i(20), ZN => n194);
   U42 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n193, ZN 
                           => n78);
   U43 : INV_X1 port map( A => i(21), ZN => n193);
   U44 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n192, ZN 
                           => n77);
   U45 : INV_X1 port map( A => i(22), ZN => n192);
   U46 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n191, ZN 
                           => n76);
   U47 : INV_X1 port map( A => i(23), ZN => n191);
   U48 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n190, ZN 
                           => n75);
   U49 : INV_X1 port map( A => i(24), ZN => n190);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n189, ZN 
                           => n74);
   U51 : INV_X1 port map( A => i(25), ZN => n189);
   U52 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n188, ZN 
                           => n73);
   U53 : INV_X1 port map( A => i(26), ZN => n188);
   U54 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n187, ZN 
                           => n72);
   U55 : INV_X1 port map( A => i(27), ZN => n187);
   U56 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n186, ZN 
                           => n71);
   U57 : INV_X1 port map( A => i(28), ZN => n186);
   U58 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U59 : INV_X1 port map( A => i(29), ZN => n185);
   U60 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U61 : INV_X1 port map( A => i(30), ZN => n184);
   U62 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U63 : INV_X1 port map( A => i(31), ZN => n183);
   U64 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U65 : INV_X1 port map( A => i(0), ZN => n214);
   U66 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U67 : INV_X1 port map( A => i(3), ZN => n211);
   U68 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U69 : INV_X1 port map( A => i(4), ZN => n210);
   U70 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U71 : INV_X1 port map( A => i(5), ZN => n209);
   U72 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U73 : INV_X1 port map( A => i(9), ZN => n205);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n216);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_7 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_7;

architecture SYN_behavioral of reg_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180, n181, n182,
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n215, Z => n177);
   U4 : BUF_X1 port map( A => n215, Z => n176);
   U5 : BUF_X1 port map( A => n215, Z => n178);
   U6 : BUF_X1 port map( A => n216, Z => n179);
   U7 : BUF_X1 port map( A => n216, Z => n180);
   U8 : BUF_X1 port map( A => n216, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n215);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n187, ZN 
                           => n99);
   U11 : INV_X1 port map( A => i(0), ZN => n187);
   U12 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n183, ZN 
                           => n95);
   U13 : INV_X1 port map( A => i(4), ZN => n183);
   U14 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n185, ZN 
                           => n97);
   U15 : INV_X1 port map( A => i(2), ZN => n185);
   U16 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n186, ZN 
                           => n98);
   U17 : INV_X1 port map( A => i(1), ZN => n186);
   U18 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n184, ZN 
                           => n96);
   U19 : INV_X1 port map( A => i(3), ZN => n184);
   U20 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n188, ZN 
                           => n94);
   U21 : INV_X1 port map( A => i(5), ZN => n188);
   U22 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n189, ZN 
                           => n93);
   U23 : INV_X1 port map( A => i(6), ZN => n189);
   U24 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n203, ZN 
                           => n79);
   U25 : INV_X1 port map( A => i(20), ZN => n203);
   U26 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n204, ZN 
                           => n78);
   U27 : INV_X1 port map( A => i(21), ZN => n204);
   U28 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n205, ZN 
                           => n77);
   U29 : INV_X1 port map( A => i(22), ZN => n205);
   U30 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n206, ZN 
                           => n76);
   U31 : INV_X1 port map( A => i(23), ZN => n206);
   U32 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n207, ZN 
                           => n75);
   U33 : INV_X1 port map( A => i(24), ZN => n207);
   U34 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n208, ZN 
                           => n74);
   U35 : INV_X1 port map( A => i(25), ZN => n208);
   U36 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n209, ZN 
                           => n73);
   U37 : INV_X1 port map( A => i(26), ZN => n209);
   U38 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n210, ZN 
                           => n72);
   U39 : INV_X1 port map( A => i(27), ZN => n210);
   U40 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n211, ZN 
                           => n71);
   U41 : INV_X1 port map( A => i(28), ZN => n211);
   U42 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n212, ZN 
                           => n70);
   U43 : INV_X1 port map( A => i(29), ZN => n212);
   U44 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n213, ZN 
                           => n69);
   U45 : INV_X1 port map( A => i(30), ZN => n213);
   U46 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n214, ZN 
                           => n68);
   U47 : INV_X1 port map( A => i(31), ZN => n214);
   U48 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n190, ZN 
                           => n92);
   U49 : INV_X1 port map( A => i(7), ZN => n190);
   U50 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n191, ZN 
                           => n91);
   U51 : INV_X1 port map( A => i(8), ZN => n191);
   U52 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n192, ZN 
                           => n90);
   U53 : INV_X1 port map( A => i(9), ZN => n192);
   U54 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n193, ZN 
                           => n89);
   U55 : INV_X1 port map( A => i(10), ZN => n193);
   U56 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n194, ZN 
                           => n88);
   U57 : INV_X1 port map( A => i(11), ZN => n194);
   U58 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n195, ZN 
                           => n87);
   U59 : INV_X1 port map( A => i(12), ZN => n195);
   U60 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n196, ZN 
                           => n86);
   U61 : INV_X1 port map( A => i(13), ZN => n196);
   U62 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n197, ZN 
                           => n85);
   U63 : INV_X1 port map( A => i(14), ZN => n197);
   U64 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n198, ZN 
                           => n84);
   U65 : INV_X1 port map( A => i(15), ZN => n198);
   U66 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n199, ZN 
                           => n83);
   U67 : INV_X1 port map( A => i(16), ZN => n199);
   U68 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n200, ZN 
                           => n82);
   U69 : INV_X1 port map( A => i(17), ZN => n200);
   U70 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n201, ZN 
                           => n81);
   U71 : INV_X1 port map( A => i(18), ZN => n201);
   U72 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n202, ZN 
                           => n80);
   U73 : INV_X1 port map( A => i(19), ZN => n202);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n216);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_4 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_4;

architecture SYN_behavioral of reg_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180, n181, n182,
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n215, Z => n177);
   U4 : BUF_X1 port map( A => n215, Z => n176);
   U5 : BUF_X1 port map( A => n215, Z => n178);
   U6 : BUF_X1 port map( A => n216, Z => n179);
   U7 : BUF_X1 port map( A => n216, Z => n180);
   U8 : BUF_X1 port map( A => n216, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n215);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U11 : INV_X1 port map( A => i(0), ZN => n214);
   U12 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U13 : INV_X1 port map( A => i(1), ZN => n213);
   U14 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U15 : INV_X1 port map( A => i(2), ZN => n212);
   U16 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U17 : INV_X1 port map( A => i(3), ZN => n211);
   U18 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U19 : INV_X1 port map( A => i(4), ZN => n210);
   U20 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U21 : INV_X1 port map( A => i(5), ZN => n209);
   U22 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U23 : INV_X1 port map( A => i(6), ZN => n208);
   U24 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U25 : INV_X1 port map( A => i(7), ZN => n207);
   U26 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U27 : INV_X1 port map( A => i(8), ZN => n206);
   U28 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U29 : INV_X1 port map( A => i(9), ZN => n205);
   U30 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U31 : INV_X1 port map( A => i(10), ZN => n204);
   U32 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U33 : INV_X1 port map( A => i(11), ZN => n203);
   U34 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U35 : INV_X1 port map( A => i(12), ZN => n202);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U37 : INV_X1 port map( A => i(13), ZN => n201);
   U38 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U39 : INV_X1 port map( A => i(14), ZN => n200);
   U40 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n199, ZN 
                           => n84);
   U41 : INV_X1 port map( A => i(15), ZN => n199);
   U42 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n198, ZN 
                           => n83);
   U43 : INV_X1 port map( A => i(16), ZN => n198);
   U44 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n197, ZN 
                           => n82);
   U45 : INV_X1 port map( A => i(17), ZN => n197);
   U46 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n196, ZN 
                           => n81);
   U47 : INV_X1 port map( A => i(18), ZN => n196);
   U48 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n195, ZN 
                           => n80);
   U49 : INV_X1 port map( A => i(19), ZN => n195);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n194, ZN 
                           => n79);
   U51 : INV_X1 port map( A => i(20), ZN => n194);
   U52 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n193, ZN 
                           => n78);
   U53 : INV_X1 port map( A => i(21), ZN => n193);
   U54 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n192, ZN 
                           => n77);
   U55 : INV_X1 port map( A => i(22), ZN => n192);
   U56 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n191, ZN 
                           => n76);
   U57 : INV_X1 port map( A => i(23), ZN => n191);
   U58 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n190, ZN 
                           => n75);
   U59 : INV_X1 port map( A => i(24), ZN => n190);
   U60 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n189, ZN 
                           => n74);
   U61 : INV_X1 port map( A => i(25), ZN => n189);
   U62 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n188, ZN 
                           => n73);
   U63 : INV_X1 port map( A => i(26), ZN => n188);
   U64 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n187, ZN 
                           => n72);
   U65 : INV_X1 port map( A => i(27), ZN => n187);
   U66 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n186, ZN 
                           => n71);
   U67 : INV_X1 port map( A => i(28), ZN => n186);
   U68 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U69 : INV_X1 port map( A => i(29), ZN => n185);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U71 : INV_X1 port map( A => i(30), ZN => n184);
   U72 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U73 : INV_X1 port map( A => i(31), ZN => n183);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n216);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_3 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_3;

architecture SYN_behavioral of reg_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180, n181, n182,
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n215, Z => n177);
   U4 : BUF_X1 port map( A => n215, Z => n176);
   U5 : BUF_X1 port map( A => n215, Z => n178);
   U6 : BUF_X1 port map( A => n216, Z => n179);
   U7 : BUF_X1 port map( A => n216, Z => n180);
   U8 : BUF_X1 port map( A => n216, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n215);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U11 : INV_X1 port map( A => i(0), ZN => n214);
   U12 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U13 : INV_X1 port map( A => i(1), ZN => n213);
   U14 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U15 : INV_X1 port map( A => i(2), ZN => n212);
   U16 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U17 : INV_X1 port map( A => i(3), ZN => n211);
   U18 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U19 : INV_X1 port map( A => i(4), ZN => n210);
   U20 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U21 : INV_X1 port map( A => i(5), ZN => n209);
   U22 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U23 : INV_X1 port map( A => i(6), ZN => n208);
   U24 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U25 : INV_X1 port map( A => i(7), ZN => n207);
   U26 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U27 : INV_X1 port map( A => i(8), ZN => n206);
   U28 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U29 : INV_X1 port map( A => i(9), ZN => n205);
   U30 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U31 : INV_X1 port map( A => i(10), ZN => n204);
   U32 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U33 : INV_X1 port map( A => i(11), ZN => n203);
   U34 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U35 : INV_X1 port map( A => i(12), ZN => n202);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U37 : INV_X1 port map( A => i(13), ZN => n201);
   U38 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U39 : INV_X1 port map( A => i(14), ZN => n200);
   U40 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n199, ZN 
                           => n84);
   U41 : INV_X1 port map( A => i(15), ZN => n199);
   U42 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n198, ZN 
                           => n83);
   U43 : INV_X1 port map( A => i(16), ZN => n198);
   U44 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n197, ZN 
                           => n82);
   U45 : INV_X1 port map( A => i(17), ZN => n197);
   U46 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n196, ZN 
                           => n81);
   U47 : INV_X1 port map( A => i(18), ZN => n196);
   U48 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n195, ZN 
                           => n80);
   U49 : INV_X1 port map( A => i(19), ZN => n195);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n194, ZN 
                           => n79);
   U51 : INV_X1 port map( A => i(20), ZN => n194);
   U52 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n193, ZN 
                           => n78);
   U53 : INV_X1 port map( A => i(21), ZN => n193);
   U54 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n192, ZN 
                           => n77);
   U55 : INV_X1 port map( A => i(22), ZN => n192);
   U56 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n191, ZN 
                           => n76);
   U57 : INV_X1 port map( A => i(23), ZN => n191);
   U58 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n190, ZN 
                           => n75);
   U59 : INV_X1 port map( A => i(24), ZN => n190);
   U60 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n189, ZN 
                           => n74);
   U61 : INV_X1 port map( A => i(25), ZN => n189);
   U62 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n188, ZN 
                           => n73);
   U63 : INV_X1 port map( A => i(26), ZN => n188);
   U64 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n187, ZN 
                           => n72);
   U65 : INV_X1 port map( A => i(27), ZN => n187);
   U66 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n186, ZN 
                           => n71);
   U67 : INV_X1 port map( A => i(28), ZN => n186);
   U68 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U69 : INV_X1 port map( A => i(29), ZN => n185);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U71 : INV_X1 port map( A => i(30), ZN => n184);
   U72 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U73 : INV_X1 port map( A => i(31), ZN => n183);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n216);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_1 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_1;

architecture SYN_behavioral of reg_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180, n181, n182,
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n215, Z => n177);
   U4 : BUF_X1 port map( A => n215, Z => n176);
   U5 : BUF_X1 port map( A => n215, Z => n178);
   U6 : BUF_X1 port map( A => n216, Z => n179);
   U7 : BUF_X1 port map( A => n216, Z => n180);
   U8 : BUF_X1 port map( A => n216, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n215);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U11 : INV_X1 port map( A => i(0), ZN => n214);
   U12 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U13 : INV_X1 port map( A => i(1), ZN => n213);
   U14 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U15 : INV_X1 port map( A => i(2), ZN => n212);
   U16 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U17 : INV_X1 port map( A => i(3), ZN => n211);
   U18 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U19 : INV_X1 port map( A => i(4), ZN => n210);
   U20 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U21 : INV_X1 port map( A => i(5), ZN => n209);
   U22 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U23 : INV_X1 port map( A => i(6), ZN => n208);
   U24 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U25 : INV_X1 port map( A => i(7), ZN => n207);
   U26 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U27 : INV_X1 port map( A => i(8), ZN => n206);
   U28 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U29 : INV_X1 port map( A => i(9), ZN => n205);
   U30 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U31 : INV_X1 port map( A => i(10), ZN => n204);
   U32 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U33 : INV_X1 port map( A => i(11), ZN => n203);
   U34 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U35 : INV_X1 port map( A => i(12), ZN => n202);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U37 : INV_X1 port map( A => i(13), ZN => n201);
   U38 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U39 : INV_X1 port map( A => i(14), ZN => n200);
   U40 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n199, ZN 
                           => n84);
   U41 : INV_X1 port map( A => i(15), ZN => n199);
   U42 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n198, ZN 
                           => n83);
   U43 : INV_X1 port map( A => i(16), ZN => n198);
   U44 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n197, ZN 
                           => n82);
   U45 : INV_X1 port map( A => i(17), ZN => n197);
   U46 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n196, ZN 
                           => n81);
   U47 : INV_X1 port map( A => i(18), ZN => n196);
   U48 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n195, ZN 
                           => n80);
   U49 : INV_X1 port map( A => i(19), ZN => n195);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n194, ZN 
                           => n79);
   U51 : INV_X1 port map( A => i(20), ZN => n194);
   U52 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n193, ZN 
                           => n78);
   U53 : INV_X1 port map( A => i(21), ZN => n193);
   U54 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n192, ZN 
                           => n77);
   U55 : INV_X1 port map( A => i(22), ZN => n192);
   U56 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n191, ZN 
                           => n76);
   U57 : INV_X1 port map( A => i(23), ZN => n191);
   U58 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n190, ZN 
                           => n75);
   U59 : INV_X1 port map( A => i(24), ZN => n190);
   U60 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n189, ZN 
                           => n74);
   U61 : INV_X1 port map( A => i(25), ZN => n189);
   U62 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n188, ZN 
                           => n73);
   U63 : INV_X1 port map( A => i(26), ZN => n188);
   U64 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n187, ZN 
                           => n72);
   U65 : INV_X1 port map( A => i(27), ZN => n187);
   U66 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n186, ZN 
                           => n71);
   U67 : INV_X1 port map( A => i(28), ZN => n186);
   U68 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U69 : INV_X1 port map( A => i(29), ZN => n185);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U71 : INV_X1 port map( A => i(30), ZN => n184);
   U72 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U73 : INV_X1 port map( A => i(31), ZN => n183);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n216);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_26 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_26;

architecture SYN_BEHAVIORAL of PG_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_25 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_25;

architecture SYN_BEHAVIORAL of PG_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_24 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_24;

architecture SYN_BEHAVIORAL of PG_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_23 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_23;

architecture SYN_BEHAVIORAL of PG_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => g_Out);
   U2 : INV_X1 port map( A => g2, ZN => n7);
   U3 : INV_X1 port map( A => p1, ZN => n8);
   U4 : INV_X1 port map( A => g1, ZN => n9);
   U5 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_22 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_22;

architecture SYN_BEHAVIORAL of PG_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U2 : INV_X1 port map( A => n8, ZN => g_Out);
   U3 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_21 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_21;

architecture SYN_BEHAVIORAL of PG_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => g_Out);
   U2 : INV_X1 port map( A => g2, ZN => n7);
   U3 : INV_X1 port map( A => p1, ZN => n8);
   U4 : INV_X1 port map( A => g1, ZN => n9);
   U5 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_20 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_20;

architecture SYN_BEHAVIORAL of PG_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_19 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_19;

architecture SYN_BEHAVIORAL of PG_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_18 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_18;

architecture SYN_BEHAVIORAL of PG_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_17 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_17;

architecture SYN_BEHAVIORAL of PG_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U2 : INV_X1 port map( A => n8, ZN => g_Out);
   U3 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_16 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_16;

architecture SYN_BEHAVIORAL of PG_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_15 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_15;

architecture SYN_BEHAVIORAL of PG_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_14 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_14;

architecture SYN_BEHAVIORAL of PG_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U2 : INV_X1 port map( A => n8, ZN => g_Out);
   U3 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_13 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_13;

architecture SYN_BEHAVIORAL of PG_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U2 : INV_X1 port map( A => n8, ZN => g_Out);
   U3 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_12 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_12;

architecture SYN_BEHAVIORAL of PG_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U2 : INV_X1 port map( A => n8, ZN => g_Out);
   U3 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_11 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_11;

architecture SYN_BEHAVIORAL of PG_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_10 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_10;

architecture SYN_BEHAVIORAL of PG_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_9 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_9;

architecture SYN_BEHAVIORAL of PG_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_8 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_8;

architecture SYN_BEHAVIORAL of PG_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_7 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_7;

architecture SYN_BEHAVIORAL of PG_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_6 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_6;

architecture SYN_BEHAVIORAL of PG_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_5 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_5;

architecture SYN_BEHAVIORAL of PG_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_4 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_4;

architecture SYN_BEHAVIORAL of PG_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U3 : INV_X1 port map( A => n8, ZN => g_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_3 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_3;

architecture SYN_BEHAVIORAL of PG_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U2 : INV_X1 port map( A => n8, ZN => g_Out);
   U3 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_2 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_2;

architecture SYN_BEHAVIORAL of PG_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U3 : INV_X1 port map( A => n8, ZN => g_Out);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_1 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_1;

architecture SYN_BEHAVIORAL of PG_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n8, ZN => g_Out);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U3 : AOI21_X1 port map( B1 => g2, B2 => p1, A => g1, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_5 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_5;

architecture SYN_behavioral of reg_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180, n181, n182,
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n215, Z => n177);
   U4 : BUF_X1 port map( A => n215, Z => n176);
   U5 : BUF_X1 port map( A => n215, Z => n178);
   U6 : BUF_X1 port map( A => n216, Z => n179);
   U7 : BUF_X1 port map( A => n216, Z => n180);
   U8 : BUF_X1 port map( A => n216, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n215);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U11 : INV_X1 port map( A => i(0), ZN => n214);
   U12 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U13 : INV_X1 port map( A => i(1), ZN => n213);
   U14 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U15 : INV_X1 port map( A => i(2), ZN => n212);
   U16 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U17 : INV_X1 port map( A => i(3), ZN => n211);
   U18 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U19 : INV_X1 port map( A => i(4), ZN => n210);
   U20 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U21 : INV_X1 port map( A => i(5), ZN => n209);
   U22 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U23 : INV_X1 port map( A => i(6), ZN => n208);
   U24 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U25 : INV_X1 port map( A => i(7), ZN => n207);
   U26 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U27 : INV_X1 port map( A => i(8), ZN => n206);
   U28 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U29 : INV_X1 port map( A => i(9), ZN => n205);
   U30 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U31 : INV_X1 port map( A => i(10), ZN => n204);
   U32 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U33 : INV_X1 port map( A => i(11), ZN => n203);
   U34 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U35 : INV_X1 port map( A => i(12), ZN => n202);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U37 : INV_X1 port map( A => i(13), ZN => n201);
   U38 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U39 : INV_X1 port map( A => i(14), ZN => n200);
   U40 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n199, ZN 
                           => n84);
   U41 : INV_X1 port map( A => i(15), ZN => n199);
   U42 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n198, ZN 
                           => n83);
   U43 : INV_X1 port map( A => i(16), ZN => n198);
   U44 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n197, ZN 
                           => n82);
   U45 : INV_X1 port map( A => i(17), ZN => n197);
   U46 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n196, ZN 
                           => n81);
   U47 : INV_X1 port map( A => i(18), ZN => n196);
   U48 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n195, ZN 
                           => n80);
   U49 : INV_X1 port map( A => i(19), ZN => n195);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n194, ZN 
                           => n79);
   U51 : INV_X1 port map( A => i(20), ZN => n194);
   U52 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n193, ZN 
                           => n78);
   U53 : INV_X1 port map( A => i(21), ZN => n193);
   U54 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n192, ZN 
                           => n77);
   U55 : INV_X1 port map( A => i(22), ZN => n192);
   U56 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n191, ZN 
                           => n76);
   U57 : INV_X1 port map( A => i(23), ZN => n191);
   U58 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n190, ZN 
                           => n75);
   U59 : INV_X1 port map( A => i(24), ZN => n190);
   U60 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n189, ZN 
                           => n74);
   U61 : INV_X1 port map( A => i(25), ZN => n189);
   U62 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n188, ZN 
                           => n73);
   U63 : INV_X1 port map( A => i(26), ZN => n188);
   U64 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n187, ZN 
                           => n72);
   U65 : INV_X1 port map( A => i(27), ZN => n187);
   U66 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n186, ZN 
                           => n71);
   U67 : INV_X1 port map( A => i(28), ZN => n186);
   U68 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U69 : INV_X1 port map( A => i(29), ZN => n185);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U71 : INV_X1 port map( A => i(30), ZN => n184);
   U72 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U73 : INV_X1 port map( A => i(31), ZN => n183);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n216);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_2 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_2;

architecture SYN_behavioral of reg_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180, n181, n182,
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n215, Z => n177);
   U4 : BUF_X1 port map( A => n215, Z => n176);
   U5 : BUF_X1 port map( A => n215, Z => n178);
   U6 : BUF_X1 port map( A => n216, Z => n179);
   U7 : BUF_X1 port map( A => n216, Z => n180);
   U8 : BUF_X1 port map( A => n216, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n215);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n204, ZN 
                           => n99);
   U11 : INV_X1 port map( A => i(0), ZN => n204);
   U12 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n209, ZN 
                           => n98);
   U13 : INV_X1 port map( A => i(1), ZN => n209);
   U14 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n203, ZN 
                           => n97);
   U15 : INV_X1 port map( A => i(2), ZN => n203);
   U16 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n207, ZN 
                           => n96);
   U17 : INV_X1 port map( A => i(3), ZN => n207);
   U18 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n202, ZN 
                           => n95);
   U19 : INV_X1 port map( A => i(4), ZN => n202);
   U20 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n201, ZN 
                           => n94);
   U21 : INV_X1 port map( A => i(5), ZN => n201);
   U22 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n200, ZN 
                           => n93);
   U23 : INV_X1 port map( A => i(6), ZN => n200);
   U24 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n199, ZN 
                           => n92);
   U25 : INV_X1 port map( A => i(7), ZN => n199);
   U26 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n198, ZN 
                           => n91);
   U27 : INV_X1 port map( A => i(8), ZN => n198);
   U28 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n210, ZN 
                           => n90);
   U29 : INV_X1 port map( A => i(9), ZN => n210);
   U30 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n197, ZN 
                           => n89);
   U31 : INV_X1 port map( A => i(10), ZN => n197);
   U32 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n196, ZN 
                           => n88);
   U33 : INV_X1 port map( A => i(11), ZN => n196);
   U34 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n214, ZN 
                           => n87);
   U35 : INV_X1 port map( A => i(12), ZN => n214);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n208, ZN 
                           => n86);
   U37 : INV_X1 port map( A => i(13), ZN => n208);
   U38 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n195, ZN 
                           => n85);
   U39 : INV_X1 port map( A => i(14), ZN => n195);
   U40 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n194, ZN 
                           => n84);
   U41 : INV_X1 port map( A => i(15), ZN => n194);
   U42 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n193, ZN 
                           => n83);
   U43 : INV_X1 port map( A => i(16), ZN => n193);
   U44 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n192, ZN 
                           => n82);
   U45 : INV_X1 port map( A => i(17), ZN => n192);
   U46 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n191, ZN 
                           => n81);
   U47 : INV_X1 port map( A => i(18), ZN => n191);
   U48 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n213, ZN 
                           => n80);
   U49 : INV_X1 port map( A => i(19), ZN => n213);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n211, ZN 
                           => n79);
   U51 : INV_X1 port map( A => i(20), ZN => n211);
   U52 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n190, ZN 
                           => n78);
   U53 : INV_X1 port map( A => i(21), ZN => n190);
   U54 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n189, ZN 
                           => n77);
   U55 : INV_X1 port map( A => i(22), ZN => n189);
   U56 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n205, ZN 
                           => n76);
   U57 : INV_X1 port map( A => i(23), ZN => n205);
   U58 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n188, ZN 
                           => n75);
   U59 : INV_X1 port map( A => i(24), ZN => n188);
   U60 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n206, ZN 
                           => n74);
   U61 : INV_X1 port map( A => i(25), ZN => n206);
   U62 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n187, ZN 
                           => n73);
   U63 : INV_X1 port map( A => i(26), ZN => n187);
   U64 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n186, ZN 
                           => n72);
   U65 : INV_X1 port map( A => i(27), ZN => n186);
   U66 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n212, ZN 
                           => n71);
   U67 : INV_X1 port map( A => i(28), ZN => n212);
   U68 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U69 : INV_X1 port map( A => i(29), ZN => n185);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U71 : INV_X1 port map( A => i(30), ZN => n184);
   U72 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U73 : INV_X1 port map( A => i(31), ZN => n183);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n216);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Mux21_3 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end Mux21_3;

architecture SYN_Behavioral of Mux21_3 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249 : 
      std_logic;

begin
   
   U1 : INV_X1 port map( A => n221, ZN => y(12));
   U2 : INV_X1 port map( A => n231, ZN => y(21));
   U3 : INV_X1 port map( A => n234, ZN => y(24));
   U4 : INV_X1 port map( A => n245, ZN => y(5));
   U5 : INV_X1 port map( A => n238, ZN => y(28));
   U6 : INV_X1 port map( A => n230, ZN => y(20));
   U7 : INV_X1 port map( A => n249, ZN => y(9));
   U8 : INV_X1 port map( A => n229, ZN => y(1));
   U9 : INV_X1 port map( A => n222, ZN => y(13));
   U10 : INV_X1 port map( A => n235, ZN => y(25));
   U11 : INV_X1 port map( A => n223, ZN => y(14));
   U12 : INV_X1 port map( A => n225, ZN => y(16));
   U13 : INV_X1 port map( A => n226, ZN => y(17));
   U14 : INV_X1 port map( A => n227, ZN => y(18));
   U15 : INV_X1 port map( A => n232, ZN => y(22));
   U16 : INV_X1 port map( A => n236, ZN => y(26));
   U17 : INV_X1 port map( A => n243, ZN => y(3));
   U18 : INV_X1 port map( A => n247, ZN => y(7));
   U19 : INV_X1 port map( A => n220, ZN => y(11));
   U20 : INV_X1 port map( A => n224, ZN => y(15));
   U21 : INV_X1 port map( A => n228, ZN => y(19));
   U22 : INV_X1 port map( A => n233, ZN => y(23));
   U23 : INV_X1 port map( A => n237, ZN => y(27));
   U24 : INV_X2 port map( A => n184, ZN => n173);
   U25 : MUX2_X1 port map( A => b(0), B => a(0), S => sel, Z => y(0));
   U26 : CLKBUF_X1 port map( A => n185, Z => n183);
   U27 : CLKBUF_X1 port map( A => n185, Z => n182);
   U28 : CLKBUF_X1 port map( A => sel, Z => n172);
   U29 : INV_X1 port map( A => n184, ZN => n174);
   U30 : BUF_X1 port map( A => n186, Z => n179);
   U31 : BUF_X1 port map( A => n186, Z => n178);
   U32 : BUF_X1 port map( A => n186, Z => n180);
   U33 : BUF_X1 port map( A => n186, Z => n181);
   U34 : BUF_X1 port map( A => n185, Z => n184);
   U35 : BUF_X1 port map( A => n186, Z => n177);
   U36 : BUF_X1 port map( A => n186, Z => n176);
   U37 : INV_X1 port map( A => n172, ZN => n185);
   U38 : INV_X1 port map( A => n172, ZN => n186);
   U39 : INV_X1 port map( A => n241, ZN => y(30));
   U40 : AOI22_X1 port map( A1 => a(30), A2 => n174, B1 => b(30), B2 => n178, 
                           ZN => n241);
   U41 : AOI22_X1 port map( A1 => a(25), A2 => n174, B1 => b(25), B2 => n179, 
                           ZN => n235);
   U42 : AOI22_X1 port map( A1 => a(1), A2 => n173, B1 => b(1), B2 => n181, ZN 
                           => n229);
   U43 : AOI22_X1 port map( A1 => a(26), A2 => n174, B1 => b(26), B2 => n179, 
                           ZN => n236);
   U44 : AOI22_X1 port map( A1 => a(22), A2 => n174, B1 => b(22), B2 => n180, 
                           ZN => n232);
   U45 : AOI22_X1 port map( A1 => a(23), A2 => n174, B1 => b(23), B2 => n180, 
                           ZN => n233);
   U46 : INV_X1 port map( A => n242, ZN => y(31));
   U47 : AOI22_X1 port map( A1 => a(13), A2 => n173, B1 => b(13), B2 => n182, 
                           ZN => n222);
   U48 : AOI22_X1 port map( A1 => a(28), A2 => n174, B1 => b(28), B2 => n178, 
                           ZN => n238);
   U49 : AOI22_X1 port map( A1 => a(18), A2 => n173, B1 => b(18), B2 => n181, 
                           ZN => n227);
   U50 : AOI22_X1 port map( A1 => a(15), A2 => n173, B1 => b(15), B2 => n182, 
                           ZN => n224);
   U51 : AOI22_X1 port map( A1 => a(19), A2 => n173, B1 => b(19), B2 => n181, 
                           ZN => n228);
   U52 : AOI22_X1 port map( A1 => a(17), A2 => n173, B1 => b(17), B2 => n181, 
                           ZN => n226);
   U53 : AOI22_X1 port map( A1 => a(24), A2 => n174, B1 => b(24), B2 => n179, 
                           ZN => n234);
   U54 : AOI22_X1 port map( A1 => a(27), A2 => n174, B1 => b(27), B2 => n179, 
                           ZN => n237);
   U55 : AOI22_X1 port map( A1 => a(14), A2 => n173, B1 => b(14), B2 => n182, 
                           ZN => n223);
   U56 : AOI22_X1 port map( A1 => a(12), A2 => n173, B1 => b(12), B2 => n183, 
                           ZN => n221);
   U57 : AOI22_X1 port map( A1 => a(11), A2 => n173, B1 => b(11), B2 => n183, 
                           ZN => n220);
   U58 : AOI22_X1 port map( A1 => a(16), A2 => n173, B1 => b(16), B2 => n182, 
                           ZN => n225);
   U59 : AOI22_X1 port map( A1 => a(2), A2 => n174, B1 => b(2), B2 => n178, ZN 
                           => n240);
   U60 : INV_X1 port map( A => n239, ZN => y(29));
   U61 : AOI22_X1 port map( A1 => a(29), A2 => n174, B1 => b(29), B2 => n178, 
                           ZN => n239);
   U62 : AOI22_X1 port map( A1 => a(21), A2 => n174, B1 => b(21), B2 => n180, 
                           ZN => n231);
   U63 : AOI22_X1 port map( A1 => a(20), A2 => n174, B1 => b(20), B2 => n180, 
                           ZN => n230);
   U64 : AOI22_X1 port map( A1 => a(10), A2 => n173, B1 => b(10), B2 => n183, 
                           ZN => n219);
   U65 : AOI22_X1 port map( A1 => a(31), A2 => n175, B1 => b(31), B2 => n177, 
                           ZN => n242);
   U66 : AOI22_X1 port map( A1 => a(5), A2 => n175, B1 => b(5), B2 => n177, ZN 
                           => n245);
   U67 : AOI22_X1 port map( A1 => n175, A2 => a(9), B1 => b(9), B2 => n176, ZN 
                           => n249);
   U68 : AOI22_X1 port map( A1 => a(3), A2 => n175, B1 => b(3), B2 => n177, ZN 
                           => n243);
   U69 : AOI22_X1 port map( A1 => a(7), A2 => n175, B1 => b(7), B2 => n176, ZN 
                           => n247);
   U70 : AOI22_X1 port map( A1 => a(8), A2 => n175, B1 => b(8), B2 => n176, ZN 
                           => n248);
   U71 : AOI22_X1 port map( A1 => a(6), A2 => n175, B1 => b(6), B2 => n176, ZN 
                           => n246);
   U72 : AOI22_X1 port map( A1 => a(4), A2 => n175, B1 => b(4), B2 => n177, ZN 
                           => n244);
   U73 : INV_X1 port map( A => n184, ZN => n175);
   U74 : INV_X2 port map( A => n219, ZN => y(10));
   U75 : INV_X2 port map( A => n248, ZN => y(8));
   U76 : INV_X2 port map( A => n246, ZN => y(6));
   U77 : INV_X2 port map( A => n244, ZN => y(4));
   U78 : INV_X2 port map( A => n240, ZN => y(2));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Mux21_2 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end Mux21_2;

architecture SYN_Behavioral of Mux21_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n43, n44, n45, net132961, net132955, net132953, net132951, net132949,
      net132947, net132943, net132941, net132937, net132935, n172, n173, n174, 
      n175, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n174, ZN => net132937);
   U2 : INV_X1 port map( A => n174, ZN => net132935);
   U3 : INV_X1 port map( A => n213, ZN => y(1));
   U4 : BUF_X1 port map( A => n175, Z => n174);
   U5 : MUX2_X1 port map( A => b(12), B => a(12), S => sel, Z => y(12));
   U6 : MUX2_X1 port map( A => b(16), B => a(16), S => sel, Z => y(16));
   U7 : MUX2_X1 port map( A => b(6), B => a(6), S => sel, Z => y(6));
   U8 : MUX2_X1 port map( A => b(24), B => a(24), S => sel, Z => y(24));
   U9 : INV_X1 port map( A => n43, ZN => y(2));
   U10 : AOI22_X1 port map( A1 => a(30), A2 => net132937, B1 => b(30), B2 => 
                           n173, ZN => n172);
   U11 : INV_X1 port map( A => n172, ZN => y(30));
   U12 : BUF_X1 port map( A => n175, Z => n173);
   U13 : AOI22_X1 port map( A1 => a(28), A2 => net132937, B1 => b(28), B2 => 
                           n173, ZN => n45);
   U14 : AOI22_X1 port map( A1 => a(2), A2 => net132937, B1 => b(2), B2 => n173
                           , ZN => n43);
   U15 : AOI22_X1 port map( A1 => a(29), A2 => net132937, B1 => b(29), B2 => 
                           n173, ZN => n44);
   U16 : CLKBUF_X1 port map( A => n175, Z => net132943);
   U17 : BUF_X1 port map( A => net132961, Z => net132941);
   U18 : INV_X1 port map( A => sel, ZN => net132961);
   U19 : INV_X1 port map( A => sel, ZN => n175);
   U20 : BUF_X1 port map( A => n175, Z => net132953);
   U21 : BUF_X1 port map( A => n175, Z => net132955);
   U22 : INV_X1 port map( A => n220, ZN => y(27));
   U23 : INV_X1 port map( A => n226, ZN => y(8));
   U24 : INV_X1 port map( A => n214, ZN => y(20));
   U25 : INV_X1 port map( A => n206, ZN => y(11));
   U26 : INV_X1 port map( A => n225, ZN => y(7));
   U27 : INV_X1 port map( A => n227, ZN => y(9));
   U28 : INV_X1 port map( A => n208, ZN => y(14));
   U29 : INV_X1 port map( A => n215, ZN => y(21));
   U30 : INV_X1 port map( A => n44, ZN => y(29));
   U31 : INV_X1 port map( A => n209, ZN => y(15));
   U32 : INV_X1 port map( A => n45, ZN => y(28));
   U33 : INV_X1 port map( A => n218, ZN => y(25));
   U34 : INV_X1 port map( A => n207, ZN => y(13));
   U35 : INV_X1 port map( A => n217, ZN => y(23));
   U36 : INV_X1 port map( A => n205, ZN => y(10));
   U37 : INV_X1 port map( A => n211, ZN => y(18));
   U38 : INV_X1 port map( A => n210, ZN => y(17));
   U39 : BUF_X1 port map( A => net132961, Z => net132949);
   U40 : BUF_X1 port map( A => net132961, Z => net132951);
   U41 : BUF_X1 port map( A => net132961, Z => net132947);
   U42 : AOI22_X1 port map( A1 => net132935, A2 => a(9), B1 => b(9), B2 => 
                           net132941, ZN => n227);
   U43 : INV_X1 port map( A => n219, ZN => y(26));
   U44 : AOI22_X1 port map( A1 => a(14), A2 => net132935, B1 => b(14), B2 => 
                           net132953, ZN => n208);
   U45 : AOI22_X1 port map( A1 => a(15), A2 => net132935, B1 => b(15), B2 => 
                           net132953, ZN => n209);
   U46 : INV_X1 port map( A => n204, ZN => y(0));
   U47 : AOI22_X1 port map( A1 => a(0), A2 => net132935, B1 => b(0), B2 => 
                           net132955, ZN => n204);
   U48 : AOI22_X1 port map( A1 => a(21), A2 => net132937, B1 => b(21), B2 => 
                           net132949, ZN => n215);
   U49 : AOI22_X1 port map( A1 => a(20), A2 => net132937, B1 => b(20), B2 => 
                           net132949, ZN => n214);
   U50 : AOI22_X1 port map( A1 => a(1), A2 => net132935, B1 => b(1), B2 => 
                           net132951, ZN => n213);
   U51 : INV_X1 port map( A => n222, ZN => y(3));
   U52 : AOI22_X1 port map( A1 => a(3), A2 => net132937, B1 => b(3), B2 => 
                           net132943, ZN => n222);
   U53 : INV_X1 port map( A => n223, ZN => y(4));
   U54 : AOI22_X1 port map( A1 => a(4), A2 => net132935, B1 => b(4), B2 => 
                           net132943, ZN => n223);
   U55 : INV_X1 port map( A => n224, ZN => y(5));
   U56 : AOI22_X1 port map( A1 => a(5), A2 => net132937, B1 => b(5), B2 => 
                           net132943, ZN => n224);
   U57 : AOI22_X1 port map( A1 => a(11), A2 => net132935, B1 => b(11), B2 => 
                           net132955, ZN => n206);
   U58 : INV_X1 port map( A => n221, ZN => y(31));
   U59 : INV_X1 port map( A => n212, ZN => y(19));
   U60 : AOI22_X1 port map( A1 => a(10), A2 => net132935, B1 => b(10), B2 => 
                           net132955, ZN => n205);
   U61 : AOI22_X1 port map( A1 => a(27), A2 => net132937, B1 => b(27), B2 => 
                           net132947, ZN => n220);
   U62 : AOI22_X1 port map( A1 => a(7), A2 => net132935, B1 => b(7), B2 => 
                           net132941, ZN => n225);
   U63 : INV_X1 port map( A => n216, ZN => y(22));
   U64 : AOI22_X1 port map( A1 => a(22), A2 => net132937, B1 => b(22), B2 => 
                           net132949, ZN => n216);
   U65 : AOI22_X1 port map( A1 => a(17), A2 => net132935, B1 => b(17), B2 => 
                           net132951, ZN => n210);
   U66 : AOI22_X1 port map( A1 => a(25), A2 => net132937, B1 => b(25), B2 => 
                           net132947, ZN => n218);
   U67 : AOI22_X1 port map( A1 => a(18), A2 => net132935, B1 => b(18), B2 => 
                           net132951, ZN => n211);
   U68 : AOI22_X1 port map( A1 => a(26), A2 => net132937, B1 => b(26), B2 => 
                           net132947, ZN => n219);
   U69 : AOI22_X1 port map( A1 => a(19), A2 => net132935, B1 => b(19), B2 => 
                           net132951, ZN => n212);
   U70 : AOI22_X1 port map( A1 => a(8), A2 => net132937, B1 => b(8), B2 => 
                           net132941, ZN => n226);
   U71 : AOI22_X1 port map( A1 => a(31), A2 => net132935, B1 => b(31), B2 => 
                           net132943, ZN => n221);
   U72 : AOI22_X1 port map( A1 => a(23), A2 => net132937, B1 => b(23), B2 => 
                           net132949, ZN => n217);
   U73 : AOI22_X1 port map( A1 => a(13), A2 => net132935, B1 => b(13), B2 => 
                           net132953, ZN => n207);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Mux21_1 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end Mux21_1;

architecture SYN_Behavioral of Mux21_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n181, ZN => n172);
   U2 : BUF_X1 port map( A => n182, Z => n173);
   U3 : BUF_X1 port map( A => n173, Z => n180);
   U4 : BUF_X1 port map( A => n175, Z => n179);
   U5 : BUF_X1 port map( A => n182, Z => n178);
   U6 : BUF_X1 port map( A => n182, Z => n177);
   U7 : BUF_X1 port map( A => n182, Z => n176);
   U8 : BUF_X1 port map( A => n182, Z => n175);
   U9 : BUF_X1 port map( A => n182, Z => n174);
   U10 : BUF_X1 port map( A => n182, Z => n181);
   U11 : INV_X1 port map( A => sel, ZN => n182);
   U12 : INV_X1 port map( A => n240, ZN => y(3));
   U13 : AOI22_X1 port map( A1 => a(3), A2 => n172, B1 => b(3), B2 => n174, ZN 
                           => n240);
   U14 : INV_X1 port map( A => n241, ZN => y(4));
   U15 : AOI22_X1 port map( A1 => a(4), A2 => n172, B1 => b(4), B2 => n174, ZN 
                           => n241);
   U16 : INV_X1 port map( A => n242, ZN => y(5));
   U17 : AOI22_X1 port map( A1 => a(5), A2 => n172, B1 => b(5), B2 => n174, ZN 
                           => n242);
   U18 : INV_X1 port map( A => n243, ZN => y(6));
   U19 : AOI22_X1 port map( A1 => a(6), A2 => n172, B1 => b(6), B2 => n173, ZN 
                           => n243);
   U20 : INV_X1 port map( A => n244, ZN => y(7));
   U21 : AOI22_X1 port map( A1 => a(7), A2 => n172, B1 => b(7), B2 => n173, ZN 
                           => n244);
   U22 : INV_X1 port map( A => n245, ZN => y(8));
   U23 : AOI22_X1 port map( A1 => a(8), A2 => n172, B1 => b(8), B2 => n173, ZN 
                           => n245);
   U24 : INV_X1 port map( A => n239, ZN => y(31));
   U25 : AOI22_X1 port map( A1 => a(31), A2 => sel, B1 => b(31), B2 => n174, ZN
                           => n239);
   U26 : INV_X1 port map( A => n215, ZN => y(0));
   U27 : AOI22_X1 port map( A1 => a(0), A2 => n172, B1 => b(0), B2 => n180, ZN 
                           => n215);
   U28 : INV_X1 port map( A => n226, ZN => y(1));
   U29 : AOI22_X1 port map( A1 => a(1), A2 => n172, B1 => b(1), B2 => n178, ZN 
                           => n226);
   U30 : INV_X1 port map( A => n237, ZN => y(2));
   U31 : AOI22_X1 port map( A1 => a(2), A2 => sel, B1 => b(2), B2 => n175, ZN 
                           => n237);
   U32 : INV_X1 port map( A => n216, ZN => y(10));
   U33 : AOI22_X1 port map( A1 => a(10), A2 => n172, B1 => b(10), B2 => n180, 
                           ZN => n216);
   U34 : INV_X1 port map( A => n217, ZN => y(11));
   U35 : AOI22_X1 port map( A1 => a(11), A2 => n172, B1 => b(11), B2 => n180, 
                           ZN => n217);
   U36 : INV_X1 port map( A => n218, ZN => y(12));
   U37 : AOI22_X1 port map( A1 => a(12), A2 => n172, B1 => b(12), B2 => n180, 
                           ZN => n218);
   U38 : INV_X1 port map( A => n219, ZN => y(13));
   U39 : AOI22_X1 port map( A1 => a(13), A2 => n172, B1 => b(13), B2 => n179, 
                           ZN => n219);
   U40 : INV_X1 port map( A => n220, ZN => y(14));
   U41 : AOI22_X1 port map( A1 => a(14), A2 => n172, B1 => b(14), B2 => n179, 
                           ZN => n220);
   U42 : INV_X1 port map( A => n221, ZN => y(15));
   U43 : AOI22_X1 port map( A1 => a(15), A2 => n172, B1 => b(15), B2 => n179, 
                           ZN => n221);
   U44 : INV_X1 port map( A => n222, ZN => y(16));
   U45 : AOI22_X1 port map( A1 => a(16), A2 => n172, B1 => b(16), B2 => n179, 
                           ZN => n222);
   U46 : INV_X1 port map( A => n223, ZN => y(17));
   U47 : AOI22_X1 port map( A1 => a(17), A2 => n172, B1 => b(17), B2 => n178, 
                           ZN => n223);
   U48 : INV_X1 port map( A => n224, ZN => y(18));
   U49 : AOI22_X1 port map( A1 => a(18), A2 => n172, B1 => b(18), B2 => n178, 
                           ZN => n224);
   U50 : INV_X1 port map( A => n225, ZN => y(19));
   U51 : AOI22_X1 port map( A1 => a(19), A2 => n172, B1 => b(19), B2 => n178, 
                           ZN => n225);
   U52 : INV_X1 port map( A => n227, ZN => y(20));
   U53 : AOI22_X1 port map( A1 => a(20), A2 => sel, B1 => b(20), B2 => n177, ZN
                           => n227);
   U54 : INV_X1 port map( A => n228, ZN => y(21));
   U55 : AOI22_X1 port map( A1 => a(21), A2 => sel, B1 => b(21), B2 => n177, ZN
                           => n228);
   U56 : INV_X1 port map( A => n229, ZN => y(22));
   U57 : AOI22_X1 port map( A1 => a(22), A2 => sel, B1 => b(22), B2 => n177, ZN
                           => n229);
   U58 : INV_X1 port map( A => n230, ZN => y(23));
   U59 : AOI22_X1 port map( A1 => a(23), A2 => sel, B1 => b(23), B2 => n177, ZN
                           => n230);
   U60 : INV_X1 port map( A => n231, ZN => y(24));
   U61 : AOI22_X1 port map( A1 => a(24), A2 => sel, B1 => b(24), B2 => n176, ZN
                           => n231);
   U62 : INV_X1 port map( A => n232, ZN => y(25));
   U63 : AOI22_X1 port map( A1 => a(25), A2 => sel, B1 => b(25), B2 => n176, ZN
                           => n232);
   U64 : INV_X1 port map( A => n233, ZN => y(26));
   U65 : AOI22_X1 port map( A1 => a(26), A2 => sel, B1 => b(26), B2 => n176, ZN
                           => n233);
   U66 : INV_X1 port map( A => n234, ZN => y(27));
   U67 : AOI22_X1 port map( A1 => a(27), A2 => sel, B1 => b(27), B2 => n176, ZN
                           => n234);
   U68 : INV_X1 port map( A => n235, ZN => y(28));
   U69 : AOI22_X1 port map( A1 => a(28), A2 => sel, B1 => b(28), B2 => n175, ZN
                           => n235);
   U70 : INV_X1 port map( A => n236, ZN => y(29));
   U71 : AOI22_X1 port map( A1 => a(29), A2 => sel, B1 => b(29), B2 => n175, ZN
                           => n236);
   U72 : INV_X1 port map( A => n238, ZN => y(30));
   U73 : AOI22_X1 port map( A1 => a(30), A2 => sel, B1 => b(30), B2 => n175, ZN
                           => n238);
   U74 : INV_X1 port map( A => n246, ZN => y(9));
   U75 : AOI22_X1 port map( A1 => sel, A2 => a(9), B1 => b(9), B2 => n173, ZN 
                           => n246);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n3, B2 => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity RCA_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_0;

architecture SYN_STRUCTURAL of RCA_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSb_7 is

   port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : out 
         std_logic_vector (3 downto 0));

end CSb_7;

architecture SYN_STRUCTURAL of CSb_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, 
      out0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, n6, n7, 
      n8, n9, n26, n_1012, n_1013 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => out0_3_port, 
                           S(2) => out0_2_port, S(1) => out0_1_port, S(0) => 
                           out0_0_port, Co => n_1012);
   RCA1 : RCA_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => out1_3_port, 
                           S(2) => out1_2_port, S(1) => out1_1_port, S(0) => 
                           out1_0_port, Co => n_1013);
   U3 : INV_X1 port map( A => n8, ZN => s(1));
   U4 : INV_X1 port map( A => n6, ZN => s(3));
   U5 : INV_X1 port map( A => n7, ZN => s(2));
   U6 : INV_X1 port map( A => n9, ZN => s(0));
   U7 : AOI22_X1 port map( A1 => out0_1_port, A2 => n26, B1 => out1_1_port, B2 
                           => ci, ZN => n8);
   U8 : AOI22_X1 port map( A1 => out0_0_port, A2 => n26, B1 => out1_0_port, B2 
                           => ci, ZN => n9);
   U9 : AOI22_X1 port map( A1 => out0_2_port, A2 => n26, B1 => out1_2_port, B2 
                           => ci, ZN => n7);
   U10 : AOI22_X1 port map( A1 => out0_3_port, A2 => n26, B1 => out1_3_port, B2
                           => ci, ZN => n6);
   U11 : INV_X1 port map( A => ci, ZN => n26);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSb_0 is

   port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : out 
         std_logic_vector (3 downto 0));

end CSb_0;

architecture SYN_STRUCTURAL of CSb_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component RCA_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out0_3_port, out0_2_port, out0_1_port, 
      out0_0_port, out1_3_port, out1_2_port, out1_1_port, out1_0_port, n6, n7, 
      n8, n9, n18, n_1014, n_1015 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic0_port, S(3) => out0_3_port, 
                           S(2) => out0_2_port, S(1) => out0_1_port, S(0) => 
                           out0_0_port, Co => n_1014);
   RCA1 : RCA_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Ci => X_Logic1_port, S(3) => out1_3_port, 
                           S(2) => out1_2_port, S(1) => out1_1_port, S(0) => 
                           out1_0_port, Co => n_1015);
   U3 : INV_X1 port map( A => n6, ZN => s(3));
   U4 : AOI22_X1 port map( A1 => out0_3_port, A2 => n18, B1 => out1_3_port, B2 
                           => ci, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => s(2));
   U6 : AOI22_X1 port map( A1 => out0_2_port, A2 => n18, B1 => out1_2_port, B2 
                           => ci, ZN => n7);
   U7 : INV_X1 port map( A => n8, ZN => s(1));
   U8 : AOI22_X1 port map( A1 => out0_1_port, A2 => n18, B1 => out1_1_port, B2 
                           => ci, ZN => n8);
   U9 : INV_X1 port map( A => n9, ZN => s(0));
   U10 : AOI22_X1 port map( A1 => out0_0_port, A2 => n18, B1 => out1_0_port, B2
                           => ci, ZN => n9);
   U11 : INV_X1 port map( A => ci, ZN => n18);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PG_0 is

   port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);

end PG_0;

architecture SYN_BEHAVIORAL of PG_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => p_Out);
   U2 : INV_X1 port map( A => n2, ZN => g_Out);
   U3 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity G_0 is

   port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);

end G_0;

architecture SYN_BEHAVIORAL of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => g_Out);
   U2 : AOI21_X1 port map( B1 => p1, B2 => g2, A => g1, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity PGnet_0 is

   port( A, B : in std_logic;  p, g : out std_logic);

end PGnet_0;

architecture SYN_BEHAVIORAL of PGnet_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => p);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => g);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity COMPARATOR_M32_DW01_cmp6_1 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end COMPARATOR_M32_DW01_cmp6_1;

architecture SYN_rpl of COMPARATOR_M32_DW01_cmp6_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17
      , n18, n19, n20, n21, n22, n23, n26, n27, n29, n30, n31, n32, n33, n34, 
      n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n55, n56, n58, n59, n60, n61, n62, n63, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n82, n83, n86, n88
      , n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n100, n101, n103, 
      n105, n106, n107, n108, n109, n110, n111, n112, n115, n116, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n141, n142, n144, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n159, n161, n162, n163, 
      n164, n165, n167, n168, n169, n172, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n193, n194, n195, n198, n200, n201, n204, n206, n207, 
      n208, n209, n210, n211, n212, n216, n218, n225, n226, n227, n228, n231, 
      n233, n234, n237, n238, n239, n240, n241, n242, n243, n244, n245, n255, 
      n256, n257, n258, n263, n264, n268, n269, n270, n271, n272, n273, n276, 
      n278, n286, n287, n288, n289, n290, n292, n293, n294, n295, n298, n300, 
      n301, n303, n305, n306, n313, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511 : std_logic;

begin
   
   U281 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => n15, ZN => n11);
   U282 : NAND3_X1 port map( A1 => n21, A2 => n22, A3 => n23, ZN => n20);
   U283 : NAND3_X1 port map( A1 => n425, A2 => n29, A3 => n418, ZN => n22);
   U284 : NAND3_X1 port map( A1 => n39, A2 => n429, A3 => n40, ZN => n43);
   U285 : NAND3_X1 port map( A1 => n40, A2 => n52, A3 => n53, ZN => n51);
   U286 : NAND3_X1 port map( A1 => n438, A2 => n58, A3 => n432, ZN => n52);
   U287 : NAND3_X1 port map( A1 => n60, A2 => n39, A3 => n61, ZN => n50);
   U288 : NAND3_X1 port map( A1 => n76, A2 => n77, A3 => n78, ZN => n75);
   U289 : NAND3_X1 port map( A1 => n97, A2 => n457, A3 => n98, ZN => n101);
   U292 : NAND3_X1 port map( A1 => n467, A2 => n460, A3 => n118, ZN => n111);
   U293 : NAND3_X1 port map( A1 => n120, A2 => n97, A3 => n121, ZN => n109);
   U294 : NAND3_X1 port map( A1 => n132, A2 => n137, A3 => n138, ZN => n123);
   U295 : NAND3_X1 port map( A1 => n478, A2 => n144, A3 => n473, ZN => n137);
   U296 : NAND3_X1 port map( A1 => n151, A2 => n152, A3 => n153, ZN => n147);
   U297 : NAND3_X1 port map( A1 => n167, A2 => n168, A3 => n169, ZN => n164);
   U298 : NAND3_X1 port map( A1 => n27, A2 => n418, A3 => n423, ZN => n167);
   U299 : NAND3_X1 port map( A1 => n183, A2 => n431, A3 => n46, ZN => n182);
   U300 : NAND3_X1 port map( A1 => n183, A2 => n46, A3 => n41, ZN => n180);
   U301 : NAND3_X1 port map( A1 => n436, A2 => n56, A3 => n432, ZN => n195);
   U304 : NAND3_X1 port map( A1 => n216, A2 => n70, A3 => n72, ZN => n211);
   U305 : NAND3_X1 port map( A1 => n218, A2 => n1, A3 => n432, ZN => n209);
   U307 : NAND3_X1 port map( A1 => n216, A2 => n444, A3 => n70, ZN => n218);
   U308 : NAND3_X1 port map( A1 => n245, A2 => n459, A3 => n105, ZN => n244);
   U309 : NAND3_X1 port map( A1 => n245, A2 => n105, A3 => n99, ZN => n242);
   U310 : NAND3_X1 port map( A1 => n464, A2 => n116, A3 => n460, ZN => n257);
   U311 : NAND3_X1 port map( A1 => n276, A2 => n136, A3 => n133, ZN => n272);
   U312 : NAND3_X1 port map( A1 => n278, A2 => n465, A3 => n460, ZN => n270);
   U313 : NAND3_X1 port map( A1 => n276, A2 => n472, A3 => n136, ZN => n278);
   U314 : NAND3_X1 port map( A1 => n286, A2 => n287, A3 => n288, ZN => n268);
   U315 : NAND3_X1 port map( A1 => n293, A2 => n294, A3 => n295, ZN => n287);
   U1 : AOI21_X1 port map( B1 => n176, B2 => n177, A => n178, ZN => n163);
   U2 : NAND4_X1 port map( A1 => n179, A2 => n180, A3 => n181, A4 => n182, ZN 
                           => n178);
   U3 : AND3_X1 port map( A1 => n193, A2 => n194, A3 => n195, ZN => n177);
   U4 : OAI21_X1 port map( B1 => n206, B2 => n207, A => n208, ZN => n176);
   U5 : AOI21_X1 port map( B1 => n238, B2 => n239, A => n240, ZN => n206);
   U6 : NAND4_X1 port map( A1 => n241, A2 => n242, A3 => n243, A4 => n244, ZN 
                           => n240);
   U7 : NAND2_X1 port map( A1 => n268, A2 => n269, ZN => n238);
   U8 : NOR2_X1 port map( A1 => n255, A2 => n256, ZN => n239);
   U9 : OAI21_X1 port map( B1 => n47, B2 => n48, A => n49, ZN => n18);
   U10 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => n48);
   U11 : NOR2_X1 port map( A1 => n50, A2 => n51, ZN => n49);
   U12 : AOI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n47);
   U13 : INV_X1 port map( A => n55, ZN => n432);
   U14 : NOR2_X1 port map( A1 => n96, A2 => n83, ZN => n243);
   U15 : NOR2_X1 port map( A1 => n38, A2 => n26, ZN => n181);
   U16 : NOR2_X1 port map( A1 => n83, A2 => n448, ZN => n79);
   U17 : INV_X1 port map( A => n26, ZN => n418);
   U18 : NOR2_X1 port map( A1 => n96, A2 => n83, ZN => n95);
   U19 : NOR2_X1 port map( A1 => n209, A2 => n210, ZN => n208);
   U20 : NAND2_X1 port map( A1 => n211, A2 => n212, ZN => n210);
   U21 : NOR2_X1 port map( A1 => n441, A2 => n435, ZN => n212);
   U22 : NOR2_X1 port map( A1 => n38, A2 => n26, ZN => n37);
   U23 : NOR2_X1 port map( A1 => n130, A2 => n115, ZN => n129);
   U24 : NOR2_X1 port map( A1 => n447, A2 => n88, ZN => n76);
   U25 : NAND2_X1 port map( A1 => n450, A2 => n445, ZN => n77);
   U26 : AOI21_X1 port map( B1 => n79, B2 => n452, A => n441, ZN => n78);
   U27 : INV_X1 port map( A => n115, ZN => n460);
   U28 : NOR2_X1 port map( A1 => n141, A2 => n154, ZN => n153);
   U29 : NOR2_X1 port map( A1 => n141, A2 => n154, ZN => n295);
   U30 : INV_X1 port map( A => n83, ZN => n445);
   U31 : INV_X1 port map( A => n141, ZN => n473);
   U32 : INV_X1 port map( A => n8, ZN => LE);
   U33 : INV_X1 port map( A => n99, ZN => n455);
   U34 : INV_X1 port map( A => n133, ZN => n469);
   U35 : INV_X1 port map( A => n41, ZN => n427);
   U36 : INV_X1 port map( A => n130, ZN => n465);
   U37 : OAI21_X1 port map( B1 => n10, B2 => n11, A => n12, ZN => n8);
   U38 : NOR2_X1 port map( A1 => n13, A2 => n3, ZN => n12);
   U39 : AOI21_X1 port map( B1 => n18, B2 => n19, A => n20, ZN => n10);
   U40 : NAND2_X1 port map( A1 => n90, A2 => n231, ZN => n83);
   U41 : NAND2_X1 port map( A1 => n150, A2 => n298, ZN => n141);
   U42 : INV_X1 port map( A => n120, ZN => n459);
   U43 : INV_X1 port map( A => n60, ZN => n431);
   U44 : NAND4_X1 port map( A1 => n105, A2 => n103, A3 => n245, A4 => n264, ZN 
                           => n255);
   U45 : NAND2_X1 port map( A1 => n32, A2 => n172, ZN => n26);
   U46 : INV_X1 port map( A => n45, ZN => n429);
   U47 : NAND2_X1 port map( A1 => n121, A2 => n264, ZN => n115);
   U48 : NOR2_X1 port map( A1 => n270, A2 => n271, ZN => n269);
   U49 : NAND2_X1 port map( A1 => n272, A2 => n273, ZN => n271);
   U50 : NOR2_X1 port map( A1 => n83, A2 => n106, ZN => n234);
   U51 : NOR2_X1 port map( A1 => n91, A2 => n92, ZN => n74);
   U52 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => n91);
   U53 : OAI21_X1 port map( B1 => n455, B2 => n94, A => n95, ZN => n92);
   U54 : NOR2_X1 port map( A1 => n33, A2 => n34, ZN => n19);
   U55 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => n33);
   U56 : OAI21_X1 port map( B1 => n427, B2 => n36, A => n37, ZN => n34);
   U57 : AND2_X1 port map( A1 => n29, A2 => n46, ZN => n42);
   U58 : NOR2_X1 port map( A1 => n141, A2 => n144, ZN => n290);
   U59 : NOR2_X1 port map( A1 => n439, A2 => n65, ZN => n63);
   U60 : INV_X1 port map( A => n70, ZN => n439);
   U61 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n58, ZN => n65);
   U62 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => n67);
   U63 : NOR2_X1 port map( A1 => n141, A2 => n292, ZN => n289);
   U64 : NAND2_X1 port map( A1 => n435, A2 => n432, ZN => n53);
   U65 : INV_X1 port map( A => n59, ZN => n438);
   U66 : AND2_X1 port map( A1 => n16, A2 => n172, ZN => n168);
   U67 : NAND2_X1 port map( A1 => n420, A2 => n418, ZN => n169);
   U68 : NAND2_X1 port map( A1 => n476, A2 => n473, ZN => n138);
   U69 : INV_X1 port map( A => n146, ZN => n478);
   U70 : NOR2_X1 port map( A1 => n125, A2 => n126, ZN => n124);
   U71 : OAI211_X1 port map( C1 => n134, C2 => n135, A => n118, B => n136, ZN 
                           => n125);
   U72 : OAI21_X1 port map( B1 => n469, B2 => n128, A => n129, ZN => n126);
   U73 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => n135);
   U74 : NOR2_X1 port map( A1 => n450, A2 => n237, ZN => n233);
   U75 : AND2_X1 port map( A1 => n31, A2 => n32, ZN => n21);
   U76 : NAND2_X1 port map( A1 => n422, A2 => n418, ZN => n23);
   U77 : NOR2_X1 port map( A1 => n448, A2 => n453, ZN => n100);
   U78 : INV_X1 port map( A => n105, ZN => n453);
   U79 : NOR2_X1 port map( A1 => n2, A2 => n71, ZN => n62);
   U80 : AND3_X1 port map( A1 => n69, A2 => n68, A3 => n72, ZN => n2);
   U81 : NAND2_X1 port map( A1 => n432, A2 => n1, ZN => n71);
   U82 : NOR2_X1 port map( A1 => n305, A2 => n306, ZN => n286);
   U83 : AOI21_X1 port map( B1 => n289, B2 => n142, A => n290, ZN => n288);
   U84 : INV_X1 port map( A => n89, ZN => n444);
   U85 : NAND2_X1 port map( A1 => n39, A2 => n183, ZN => n41);
   U86 : NAND2_X1 port map( A1 => n146, A2 => n292, ZN => n154);
   U87 : NAND2_X1 port map( A1 => n97, A2 => n245, ZN => n99);
   U88 : NAND2_X1 port map( A1 => n82, A2 => n237, ZN => n96);
   U89 : NOR2_X1 port map( A1 => n9, A2 => n8, ZN => EQ);
   U90 : NAND2_X1 port map( A1 => n131, A2 => n276, ZN => n133);
   U91 : NAND2_X1 port map( A1 => n30, A2 => n175, ZN => n38);
   U92 : NAND2_X1 port map( A1 => n119, A2 => n263, ZN => n130);
   U93 : NAND2_X1 port map( A1 => n61, A2 => n204, ZN => n55);
   U94 : INV_X1 port map( A => n68, ZN => n441);
   U95 : NAND2_X1 port map( A1 => n69, A2 => n216, ZN => n72);
   U96 : NAND2_X1 port map( A1 => n89, A2 => n69, ZN => n88);
   U97 : INV_X1 port map( A => n198, ZN => n436);
   U98 : NOR2_X1 port map( A1 => n200, A2 => n201, ZN => n193);
   U99 : NAND2_X1 port map( A1 => n183, A2 => n204, ZN => n200);
   U100 : NAND2_X1 port map( A1 => n46, A2 => n45, ZN => n201);
   U101 : NAND2_X1 port map( A1 => n70, A2 => n66, ZN => n228);
   U102 : INV_X1 port map( A => n56, ZN => n435);
   U103 : INV_X1 port map( A => n86, ZN => n450);
   U104 : NAND2_X1 port map( A1 => n131, A2 => n132, ZN => n128);
   U105 : INV_X1 port map( A => n106, ZN => n448);
   U106 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => n36);
   U107 : NAND2_X1 port map( A1 => n97, A2 => n98, ZN => n94);
   U108 : NAND2_X1 port map( A1 => n276, A2 => n298, ZN => n305);
   U109 : NAND2_X1 port map( A1 => n136, A2 => n134, ZN => n306);
   U110 : AND2_X1 port map( A1 => n59, A2 => n198, ZN => n1);
   U111 : INV_X1 port map( A => n82, ZN => n452);
   U112 : NAND2_X1 port map( A1 => n257, A2 => n258, ZN => n256);
   U113 : NAND2_X1 port map( A1 => n462, A2 => n460, ZN => n258);
   U114 : INV_X1 port map( A => n263, ZN => n464);
   U115 : NAND2_X1 port map( A1 => n111, A2 => n112, ZN => n110);
   U116 : AND2_X1 port map( A1 => n313, A2 => n98, ZN => n112);
   U117 : OR2_X1 port map( A1 => n115, A2 => n116, ZN => n313);
   U118 : NAND2_X1 port map( A1 => n225, A2 => n226, ZN => n207);
   U119 : NOR2_X1 port map( A1 => n227, A2 => n228, ZN => n226);
   U120 : AOI21_X1 port map( B1 => n233, B2 => n445, A => n234, ZN => n225);
   U121 : NAND2_X1 port map( A1 => n216, A2 => n231, ZN => n227);
   U122 : INV_X1 port map( A => n27, ZN => n422);
   U123 : INV_X1 port map( A => n118, ZN => n462);
   U124 : INV_X1 port map( A => n90, ZN => n447);
   U125 : INV_X1 port map( A => n142, ZN => n476);
   U126 : NAND2_X1 port map( A1 => n107, A2 => n108, ZN => n73);
   U127 : NOR2_X1 port map( A1 => n109, A2 => n110, ZN => n108);
   U128 : OAI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n107);
   U129 : NAND2_X1 port map( A1 => n147, A2 => n148, ZN => n122);
   U130 : AND2_X1 port map( A1 => n150, A2 => n6, ZN => n148);
   U131 : AND2_X1 port map( A1 => n149, A2 => n131, ZN => n6);
   U132 : AND2_X1 port map( A1 => n5, A2 => n15, ZN => n165);
   U133 : AND2_X1 port map( A1 => n31, A2 => n17, ZN => n5);
   U134 : AND2_X1 port map( A1 => n132, A2 => n116, ZN => n273);
   U135 : AND2_X1 port map( A1 => n40, A2 => n27, ZN => n179);
   U136 : AND2_X1 port map( A1 => n98, A2 => n86, ZN => n241);
   U137 : INV_X1 port map( A => n30, ZN => n425);
   U138 : INV_X1 port map( A => n119, ZN => n467);
   U139 : INV_X1 port map( A => n29, ZN => n420);
   U140 : OR2_X1 port map( A1 => n58, A2 => n55, ZN => n194);
   U141 : INV_X1 port map( A => n149, ZN => n472);
   U142 : INV_X1 port map( A => n9, ZN => GE);
   U143 : INV_X1 port map( A => n103, ZN => n457);
   U144 : INV_X1 port map( A => n175, ZN => n423);
   U145 : INV_X1 port map( A => A(6), ZN => n470);
   U146 : INV_X1 port map( A => A(24), ZN => n428);
   U147 : INV_X1 port map( A => A(25), ZN => n426);
   U148 : NAND2_X1 port map( A1 => A(18), A2 => n493, ZN => n69);
   U149 : NAND2_X1 port map( A1 => A(6), A2 => n505, ZN => n131);
   U150 : NAND2_X1 port map( A1 => A(7), A2 => n504, ZN => n132);
   U151 : NAND2_X1 port map( A1 => A(12), A2 => n499, ZN => n97);
   U152 : NAND2_X1 port map( A1 => A(24), A2 => n487, ZN => n39);
   U153 : NAND2_X1 port map( A1 => A(25), A2 => n486, ZN => n40);
   U154 : INV_X1 port map( A => A(21), ZN => n434);
   U155 : NAND2_X1 port map( A1 => A(13), A2 => n498, ZN => n98);
   U156 : INV_X1 port map( A => A(22), ZN => n433);
   U157 : INV_X1 port map( A => B(2), ZN => n509);
   U158 : INV_X1 port map( A => A(14), ZN => n451);
   U159 : INV_X1 port map( A => A(23), ZN => n430);
   U160 : NAND2_X1 port map( A1 => A(19), A2 => n492, ZN => n68);
   U161 : NAND2_X1 port map( A1 => A(27), A2 => n484, ZN => n27);
   U162 : INV_X1 port map( A => B(27), ZN => n484);
   U163 : NAND2_X1 port map( A1 => A(3), A2 => n508, ZN => n142);
   U164 : INV_X1 port map( A => B(3), ZN => n508);
   U165 : NAND2_X1 port map( A1 => A(26), A2 => n485, ZN => n30);
   U166 : INV_X1 port map( A => B(26), ZN => n485);
   U167 : NAND2_X1 port map( A1 => A(8), A2 => n503, ZN => n119);
   U168 : INV_X1 port map( A => B(8), ZN => n503);
   U169 : NAND2_X1 port map( A1 => A(14), A2 => n497, ZN => n82);
   U170 : NAND2_X1 port map( A1 => A(17), A2 => n494, ZN => n89);
   U171 : INV_X1 port map( A => B(17), ZN => n494);
   U172 : INV_X1 port map( A => B(4), ZN => n507);
   U173 : NAND2_X1 port map( A1 => A(16), A2 => n495, ZN => n90);
   U174 : INV_X1 port map( A => A(28), ZN => n419);
   U175 : NAND2_X1 port map( A1 => A(23), A2 => n488, ZN => n60);
   U176 : NAND2_X1 port map( A1 => A(9), A2 => n502, ZN => n116);
   U177 : NAND2_X1 port map( A1 => A(22), A2 => n489, ZN => n61);
   U178 : NAND2_X1 port map( A1 => n161, A2 => n162, ZN => n9);
   U179 : NOR2_X1 port map( A1 => n4, A2 => n7, ZN => n161);
   U180 : OAI21_X1 port map( B1 => n163, B2 => n164, A => n165, ZN => n162);
   U181 : NAND2_X1 port map( A1 => A(15), A2 => n496, ZN => n86);
   U182 : NAND2_X1 port map( A1 => A(21), A2 => n490, ZN => n56);
   U183 : NAND2_X1 port map( A1 => A(28), A2 => n483, ZN => n32);
   U184 : NAND2_X1 port map( A1 => A(11), A2 => n500, ZN => n120);
   U185 : NAND2_X1 port map( A1 => A(20), A2 => n491, ZN => n59);
   U186 : NAND2_X1 port map( A1 => A(5), A2 => n506, ZN => n149);
   U187 : INV_X1 port map( A => B(5), ZN => n506);
   U188 : NAND2_X1 port map( A1 => A(29), A2 => n482, ZN => n31);
   U189 : INV_X1 port map( A => A(1), ZN => n479);
   U190 : INV_X1 port map( A => A(30), ZN => n416);
   U191 : INV_X1 port map( A => A(29), ZN => n417);
   U192 : NAND2_X1 port map( A1 => B(27), A2 => n421, ZN => n29);
   U193 : INV_X1 port map( A => A(27), ZN => n421);
   U194 : NAND2_X1 port map( A1 => B(4), A2 => n474, ZN => n298);
   U195 : NAND2_X1 port map( A1 => B(2), A2 => n477, ZN => n292);
   U196 : NAND2_X1 port map( A1 => B(26), A2 => n424, ZN => n175);
   U197 : INV_X1 port map( A => A(26), ZN => n424);
   U198 : NAND2_X1 port map( A1 => B(17), A2 => n443, ZN => n66);
   U199 : INV_X1 port map( A => A(17), ZN => n443);
   U200 : NAND2_X1 port map( A1 => B(8), A2 => n466, ZN => n263);
   U201 : INV_X1 port map( A => A(8), ZN => n466);
   U202 : NAND2_X1 port map( A1 => B(5), A2 => n471, ZN => n134);
   U203 : INV_X1 port map( A => A(5), ZN => n471);
   U204 : INV_X1 port map( A => A(31), ZN => n415);
   U205 : NAND2_X1 port map( A1 => B(3), A2 => n475, ZN => n144);
   U206 : INV_X1 port map( A => A(3), ZN => n475);
   U207 : INV_X1 port map( A => A(13), ZN => n454);
   U208 : INV_X1 port map( A => A(18), ZN => n442);
   U209 : INV_X1 port map( A => A(15), ZN => n449);
   U210 : INV_X1 port map( A => A(12), ZN => n456);
   U211 : INV_X1 port map( A => A(7), ZN => n468);
   U212 : INV_X1 port map( A => A(19), ZN => n440);
   U213 : INV_X1 port map( A => A(9), ZN => n463);
   U214 : INV_X1 port map( A => A(11), ZN => n458);
   U215 : INV_X1 port map( A => B(1), ZN => n510);
   U216 : AND3_X1 port map( A1 => A(30), A2 => n481, A3 => n15, ZN => n3);
   U217 : INV_X1 port map( A => A(16), ZN => n446);
   U218 : INV_X1 port map( A => A(20), ZN => n437);
   U219 : NAND2_X1 port map( A1 => n155, A2 => n156, ZN => n152);
   U220 : NAND2_X1 port map( A1 => A(0), A2 => n511, ZN => n156);
   U221 : NAND2_X1 port map( A1 => A(1), A2 => n510, ZN => n155);
   U222 : NAND2_X1 port map( A1 => n300, A2 => n301, ZN => n294);
   U223 : NAND2_X1 port map( A1 => B(1), A2 => n479, ZN => n300);
   U224 : INV_X1 port map( A => A(0), ZN => n480);
   U225 : AND2_X1 port map( A1 => n303, A2 => n142, ZN => n293);
   U226 : NAND2_X1 port map( A1 => A(1), A2 => n510, ZN => n303);
   U227 : AND2_X1 port map( A1 => n159, A2 => n144, ZN => n151);
   U228 : NAND2_X1 port map( A1 => B(1), A2 => n479, ZN => n159);
   U229 : NAND2_X1 port map( A1 => A(2), A2 => n509, ZN => n146);
   U230 : INV_X1 port map( A => A(2), ZN => n477);
   U231 : NAND2_X1 port map( A1 => A(4), A2 => n507, ZN => n150);
   U232 : INV_X1 port map( A => A(4), ZN => n474);
   U233 : NAND2_X1 port map( A1 => A(10), A2 => n501, ZN => n121);
   U234 : INV_X1 port map( A => A(10), ZN => n461);
   U235 : NAND2_X1 port map( A1 => B(14), A2 => n451, ZN => n237);
   U236 : INV_X1 port map( A => B(14), ZN => n497);
   U237 : NAND2_X1 port map( A1 => B(13), A2 => n454, ZN => n105);
   U238 : INV_X1 port map( A => B(13), ZN => n498);
   U239 : NAND2_X1 port map( A1 => B(12), A2 => n456, ZN => n245);
   U240 : INV_X1 port map( A => B(12), ZN => n499);
   U241 : AND3_X1 port map( A1 => B(30), A2 => n416, A3 => n15, ZN => n7);
   U242 : INV_X1 port map( A => B(30), ZN => n481);
   U243 : XNOR2_X1 port map( A => B(30), B => A(30), ZN => n17);
   U244 : NAND2_X1 port map( A1 => B(29), A2 => n417, ZN => n16);
   U245 : INV_X1 port map( A => B(29), ZN => n482);
   U246 : NAND2_X1 port map( A1 => B(18), A2 => n442, ZN => n216);
   U247 : INV_X1 port map( A => B(18), ZN => n493);
   U248 : NAND2_X1 port map( A1 => B(9), A2 => n463, ZN => n118);
   U249 : INV_X1 port map( A => B(9), ZN => n502);
   U250 : NAND2_X1 port map( A1 => B(19), A2 => n440, ZN => n70);
   U251 : INV_X1 port map( A => B(19), ZN => n492);
   U252 : AND2_X1 port map( A1 => B(31), A2 => n415, ZN => n4);
   U253 : NOR2_X1 port map( A1 => B(31), A2 => n415, ZN => n13);
   U254 : XNOR2_X1 port map( A => B(31), B => A(31), ZN => n15);
   U255 : NAND2_X1 port map( A1 => B(7), A2 => n468, ZN => n136);
   U256 : INV_X1 port map( A => B(7), ZN => n504);
   U257 : NAND2_X1 port map( A1 => B(21), A2 => n434, ZN => n58);
   U258 : INV_X1 port map( A => B(21), ZN => n490);
   U259 : NAND2_X1 port map( A1 => B(15), A2 => n449, ZN => n106);
   U260 : INV_X1 port map( A => B(15), ZN => n496);
   U261 : NAND2_X1 port map( A1 => B(0), A2 => n480, ZN => n301);
   U262 : INV_X1 port map( A => B(0), ZN => n511);
   U263 : NAND2_X1 port map( A1 => B(16), A2 => n446, ZN => n231);
   U264 : INV_X1 port map( A => B(16), ZN => n495);
   U265 : NAND2_X1 port map( A1 => B(20), A2 => n437, ZN => n198);
   U266 : INV_X1 port map( A => B(20), ZN => n491);
   U267 : INV_X1 port map( A => B(25), ZN => n486);
   U268 : NAND2_X1 port map( A1 => B(25), A2 => n426, ZN => n46);
   U269 : NAND2_X1 port map( A1 => B(11), A2 => n458, ZN => n103);
   U270 : INV_X1 port map( A => B(11), ZN => n500);
   U271 : NAND2_X1 port map( A1 => B(23), A2 => n430, ZN => n45);
   U272 : INV_X1 port map( A => B(23), ZN => n488);
   U273 : NAND2_X1 port map( A1 => B(24), A2 => n428, ZN => n183);
   U274 : INV_X1 port map( A => B(24), ZN => n487);
   U275 : NAND2_X1 port map( A1 => B(10), A2 => n461, ZN => n264);
   U276 : INV_X1 port map( A => B(10), ZN => n501);
   U277 : NAND2_X1 port map( A1 => B(6), A2 => n470, ZN => n276);
   U278 : INV_X1 port map( A => B(6), ZN => n505);
   U279 : NAND2_X1 port map( A1 => B(28), A2 => n419, ZN => n172);
   U280 : INV_X1 port map( A => B(28), ZN => n483);
   U290 : NAND2_X1 port map( A1 => B(22), A2 => n433, ZN => n204);
   U291 : INV_X1 port map( A => B(22), ZN => n489);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity CSA is

   port( A, B : in std_logic_vector (31 downto 0);  c : in std_logic_vector (7 
         downto 0);  s : out std_logic_vector (31 downto 0));

end CSA;

architecture SYN_STRUCTURAL of CSA is

   component CSb_1
      port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSb_2
      port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSb_3
      port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSb_4
      port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSb_5
      port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSb_6
      port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSb_7
      port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSb_0
      port( A, B : in std_logic_vector (3 downto 0);  ci : in std_logic;  s : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSbi_0 : CSb_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) => 
                           A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), ci => c(0), s(3) => s(3), s(2) => s(2), 
                           s(1) => s(1), s(0) => s(0));
   CSbi_1 : CSb_7 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5), A(0) => 
                           A(4), B(3) => B(7), B(2) => B(6), B(1) => B(5), B(0)
                           => B(4), ci => c(1), s(3) => s(7), s(2) => s(6), 
                           s(1) => s(5), s(0) => s(4));
   CSbi_2 : CSb_6 port map( A(3) => A(11), A(2) => A(10), A(1) => A(9), A(0) =>
                           A(8), B(3) => B(11), B(2) => B(10), B(1) => B(9), 
                           B(0) => B(8), ci => c(2), s(3) => s(11), s(2) => 
                           s(10), s(1) => s(9), s(0) => s(8));
   CSbi_3 : CSb_5 port map( A(3) => A(15), A(2) => A(14), A(1) => A(13), A(0) 
                           => A(12), B(3) => B(15), B(2) => B(14), B(1) => 
                           B(13), B(0) => B(12), ci => c(3), s(3) => s(15), 
                           s(2) => s(14), s(1) => s(13), s(0) => s(12));
   CSbi_4 : CSb_4 port map( A(3) => A(19), A(2) => A(18), A(1) => A(17), A(0) 
                           => A(16), B(3) => B(19), B(2) => B(18), B(1) => 
                           B(17), B(0) => B(16), ci => c(4), s(3) => s(19), 
                           s(2) => s(18), s(1) => s(17), s(0) => s(16));
   CSbi_5 : CSb_3 port map( A(3) => A(23), A(2) => A(22), A(1) => A(21), A(0) 
                           => A(20), B(3) => B(23), B(2) => B(22), B(1) => 
                           B(21), B(0) => B(20), ci => c(5), s(3) => s(23), 
                           s(2) => s(22), s(1) => s(21), s(0) => s(20));
   CSbi_6 : CSb_2 port map( A(3) => A(27), A(2) => A(26), A(1) => A(25), A(0) 
                           => A(24), B(3) => B(27), B(2) => B(26), B(1) => 
                           B(25), B(0) => B(24), ci => c(6), s(3) => s(27), 
                           s(2) => s(26), s(1) => s(25), s(0) => s(24));
   CSbi_7 : CSb_1 port map( A(3) => A(31), A(2) => A(30), A(1) => A(29), A(0) 
                           => A(28), B(3) => B(31), B(2) => B(30), B(1) => 
                           B(29), B(0) => B(28), ci => c(7), s(3) => s(31), 
                           s(2) => s(30), s(1) => s(29), s(0) => s(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Cg is

   port( A, B : in std_logic_vector (31 downto 0);  cin0 : in std_logic;  cout 
         : out std_logic_vector (7 downto 0));

end Cg;

architecture SYN_STRUCTURAL of Cg is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_1
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component G_2
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component G_3
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component G_4
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component PG_1
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_2
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component G_5
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component G_6
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component PG_3
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_4
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_5
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component G_7
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component PG_6
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_7
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_8
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_9
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_10
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_11
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_12
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component G_8
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component PG_13
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_14
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_15
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_16
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_17
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_18
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_19
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_20
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_21
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_22
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_23
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_24
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_25
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_26
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component PG_0
      port( p1, g1, p2, g2 : in std_logic;  p_Out, g_Out : out std_logic);
   end component;
   
   component G_9
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component G_0
      port( p1, g1, g2 : in std_logic;  g_Out : out std_logic);
   end component;
   
   component PGnet_1
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_2
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_3
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_4
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_5
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_6
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_7
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_8
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_9
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_10
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_11
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_12
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_13
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_14
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_15
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_16
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_17
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_18
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_19
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_20
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_21
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_22
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_23
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_24
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_25
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_26
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_27
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_28
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_29
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_30
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component PGnet_0
      port( A, B : in std_logic;  p, g : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, n3, cout_2_port, 
      n6, n7, p0, g0, gsignal_4_31_port, gsignal_4_27_port, gsignal_3_31_port, 
      gsignal_3_23_port, gsignal_3_15_port, gsignal_2_31_port, 
      gsignal_2_27_port, gsignal_2_23_port, gsignal_2_19_port, 
      gsignal_2_15_port, gsignal_2_11_port, gsignal_2_7_port, gsignal_1_31_port
      , gsignal_1_29_port, gsignal_1_27_port, gsignal_1_25_port, 
      gsignal_1_23_port, gsignal_1_21_port, gsignal_1_19_port, 
      gsignal_1_17_port, gsignal_1_15_port, gsignal_1_13_port, 
      gsignal_1_11_port, gsignal_1_9_port, gsignal_1_7_port, gsignal_1_5_port, 
      gsignal_1_3_port, gsignal_1_1_port, gsignal_0_31_port, gsignal_0_30_port,
      gsignal_0_29_port, gsignal_0_28_port, gsignal_0_27_port, 
      gsignal_0_26_port, gsignal_0_25_port, gsignal_0_24_port, 
      gsignal_0_23_port, gsignal_0_22_port, gsignal_0_21_port, 
      gsignal_0_20_port, gsignal_0_19_port, gsignal_0_18_port, 
      gsignal_0_17_port, gsignal_0_16_port, gsignal_0_15_port, 
      gsignal_0_14_port, gsignal_0_13_port, gsignal_0_12_port, 
      gsignal_0_11_port, gsignal_0_10_port, gsignal_0_9_port, gsignal_0_8_port,
      gsignal_0_7_port, gsignal_0_6_port, gsignal_0_5_port, gsignal_0_4_port, 
      gsignal_0_3_port, gsignal_0_2_port, gsignal_0_1_port, gsignal_0_0_port, 
      psignal_4_31_port, psignal_4_27_port, psignal_3_31_port, 
      psignal_3_23_port, psignal_3_15_port, psignal_2_31_port, 
      psignal_2_27_port, psignal_2_23_port, psignal_2_19_port, 
      psignal_2_15_port, psignal_2_11_port, psignal_2_7_port, psignal_1_31_port
      , psignal_1_29_port, psignal_1_27_port, psignal_1_25_port, 
      psignal_1_23_port, psignal_1_21_port, psignal_1_19_port, 
      psignal_1_17_port, psignal_1_15_port, psignal_1_13_port, 
      psignal_1_11_port, psignal_1_9_port, psignal_1_7_port, psignal_1_5_port, 
      psignal_1_3_port, psignal_0_31_port, psignal_0_30_port, psignal_0_29_port
      , psignal_0_28_port, psignal_0_27_port, psignal_0_26_port, 
      psignal_0_25_port, psignal_0_24_port, psignal_0_23_port, 
      psignal_0_22_port, psignal_0_21_port, psignal_0_20_port, 
      psignal_0_19_port, psignal_0_18_port, psignal_0_17_port, 
      psignal_0_16_port, psignal_0_15_port, psignal_0_14_port, 
      psignal_0_13_port, psignal_0_12_port, psignal_0_11_port, 
      psignal_0_10_port, psignal_0_9_port, psignal_0_8_port, psignal_0_7_port, 
      psignal_0_6_port, psignal_0_5_port, psignal_0_4_port, psignal_0_3_port, 
      psignal_0_2_port, psignal_0_1_port, cout_0_port, cout_1_port : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, n3, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => p0);
   PGN1_31 : PGnet_0 port map( A => A(31), B => B(31), p => psignal_0_31_port, 
                           g => gsignal_0_31_port);
   PGN1_30 : PGnet_30 port map( A => A(30), B => B(30), p => psignal_0_30_port,
                           g => gsignal_0_30_port);
   PGN1_29 : PGnet_29 port map( A => A(29), B => B(29), p => psignal_0_29_port,
                           g => gsignal_0_29_port);
   PGN1_28 : PGnet_28 port map( A => A(28), B => B(28), p => psignal_0_28_port,
                           g => gsignal_0_28_port);
   PGN1_27 : PGnet_27 port map( A => A(27), B => B(27), p => psignal_0_27_port,
                           g => gsignal_0_27_port);
   PGN1_26 : PGnet_26 port map( A => A(26), B => B(26), p => psignal_0_26_port,
                           g => gsignal_0_26_port);
   PGN1_25 : PGnet_25 port map( A => A(25), B => B(25), p => psignal_0_25_port,
                           g => gsignal_0_25_port);
   PGN1_24 : PGnet_24 port map( A => A(24), B => B(24), p => psignal_0_24_port,
                           g => gsignal_0_24_port);
   PGN1_23 : PGnet_23 port map( A => A(23), B => B(23), p => psignal_0_23_port,
                           g => gsignal_0_23_port);
   PGN1_22 : PGnet_22 port map( A => A(22), B => B(22), p => psignal_0_22_port,
                           g => gsignal_0_22_port);
   PGN1_21 : PGnet_21 port map( A => A(21), B => B(21), p => psignal_0_21_port,
                           g => gsignal_0_21_port);
   PGN1_20 : PGnet_20 port map( A => A(20), B => B(20), p => psignal_0_20_port,
                           g => gsignal_0_20_port);
   PGN1_19 : PGnet_19 port map( A => A(19), B => B(19), p => psignal_0_19_port,
                           g => gsignal_0_19_port);
   PGN1_18 : PGnet_18 port map( A => A(18), B => B(18), p => psignal_0_18_port,
                           g => gsignal_0_18_port);
   PGN1_17 : PGnet_17 port map( A => A(17), B => B(17), p => psignal_0_17_port,
                           g => gsignal_0_17_port);
   PGN1_16 : PGnet_16 port map( A => A(16), B => B(16), p => psignal_0_16_port,
                           g => gsignal_0_16_port);
   PGN1_15 : PGnet_15 port map( A => A(15), B => B(15), p => psignal_0_15_port,
                           g => gsignal_0_15_port);
   PGN1_14 : PGnet_14 port map( A => A(14), B => B(14), p => psignal_0_14_port,
                           g => gsignal_0_14_port);
   PGN1_13 : PGnet_13 port map( A => A(13), B => B(13), p => psignal_0_13_port,
                           g => gsignal_0_13_port);
   PGN1_12 : PGnet_12 port map( A => A(12), B => B(12), p => psignal_0_12_port,
                           g => gsignal_0_12_port);
   PGN1_11 : PGnet_11 port map( A => A(11), B => B(11), p => psignal_0_11_port,
                           g => gsignal_0_11_port);
   PGN1_10 : PGnet_10 port map( A => A(10), B => B(10), p => psignal_0_10_port,
                           g => gsignal_0_10_port);
   PGN1_9 : PGnet_9 port map( A => A(9), B => B(9), p => psignal_0_9_port, g =>
                           gsignal_0_9_port);
   PGN1_8 : PGnet_8 port map( A => A(8), B => B(8), p => psignal_0_8_port, g =>
                           gsignal_0_8_port);
   PGN1_7 : PGnet_7 port map( A => A(7), B => B(7), p => psignal_0_7_port, g =>
                           gsignal_0_7_port);
   PGN1_6 : PGnet_6 port map( A => A(6), B => B(6), p => psignal_0_6_port, g =>
                           gsignal_0_6_port);
   PGN1_5 : PGnet_5 port map( A => A(5), B => B(5), p => psignal_0_5_port, g =>
                           gsignal_0_5_port);
   PGN1_4 : PGnet_4 port map( A => A(4), B => B(4), p => psignal_0_4_port, g =>
                           gsignal_0_4_port);
   PGN1_3 : PGnet_3 port map( A => A(3), B => B(3), p => psignal_0_3_port, g =>
                           gsignal_0_3_port);
   PGN1_2 : PGnet_2 port map( A => A(2), B => B(2), p => psignal_0_2_port, g =>
                           gsignal_0_2_port);
   PGN1_1 : PGnet_1 port map( A => A(1), B => B(1), p => psignal_0_1_port, g =>
                           gsignal_0_1_port);
   PGN0_0 : G_0 port map( p1 => p0, g1 => g0, g2 => cin0, g_Out => 
                           gsignal_0_0_port);
   g0_0_1 : G_9 port map( p1 => psignal_0_1_port, g1 => gsignal_0_1_port, g2 =>
                           gsignal_0_0_port, g_Out => gsignal_1_1_port);
   PGelements_0_3 : PG_0 port map( p1 => psignal_0_3_port, g1 => 
                           gsignal_0_3_port, p2 => psignal_0_2_port, g2 => 
                           gsignal_0_2_port, p_Out => psignal_1_3_port, g_Out 
                           => gsignal_1_3_port);
   PGelements_0_5 : PG_26 port map( p1 => psignal_0_5_port, g1 => 
                           gsignal_0_5_port, p2 => psignal_0_4_port, g2 => 
                           gsignal_0_4_port, p_Out => psignal_1_5_port, g_Out 
                           => gsignal_1_5_port);
   PGelements_0_7 : PG_25 port map( p1 => psignal_0_7_port, g1 => 
                           gsignal_0_7_port, p2 => psignal_0_6_port, g2 => 
                           gsignal_0_6_port, p_Out => psignal_1_7_port, g_Out 
                           => gsignal_1_7_port);
   PGelements_0_9 : PG_24 port map( p1 => psignal_0_9_port, g1 => 
                           gsignal_0_9_port, p2 => psignal_0_8_port, g2 => 
                           gsignal_0_8_port, p_Out => psignal_1_9_port, g_Out 
                           => gsignal_1_9_port);
   PGelements_0_11 : PG_23 port map( p1 => psignal_0_11_port, g1 => 
                           gsignal_0_11_port, p2 => psignal_0_10_port, g2 => 
                           gsignal_0_10_port, p_Out => psignal_1_11_port, g_Out
                           => gsignal_1_11_port);
   PGelements_0_13 : PG_22 port map( p1 => psignal_0_13_port, g1 => 
                           gsignal_0_13_port, p2 => psignal_0_12_port, g2 => 
                           gsignal_0_12_port, p_Out => psignal_1_13_port, g_Out
                           => gsignal_1_13_port);
   PGelements_0_15 : PG_21 port map( p1 => psignal_0_15_port, g1 => 
                           gsignal_0_15_port, p2 => psignal_0_14_port, g2 => 
                           gsignal_0_14_port, p_Out => psignal_1_15_port, g_Out
                           => gsignal_1_15_port);
   PGelements_0_17 : PG_20 port map( p1 => psignal_0_17_port, g1 => 
                           gsignal_0_17_port, p2 => psignal_0_16_port, g2 => 
                           gsignal_0_16_port, p_Out => psignal_1_17_port, g_Out
                           => gsignal_1_17_port);
   PGelements_0_19 : PG_19 port map( p1 => psignal_0_19_port, g1 => 
                           gsignal_0_19_port, p2 => psignal_0_18_port, g2 => 
                           gsignal_0_18_port, p_Out => psignal_1_19_port, g_Out
                           => gsignal_1_19_port);
   PGelements_0_21 : PG_18 port map( p1 => psignal_0_21_port, g1 => 
                           gsignal_0_21_port, p2 => psignal_0_20_port, g2 => 
                           gsignal_0_20_port, p_Out => psignal_1_21_port, g_Out
                           => gsignal_1_21_port);
   PGelements_0_23 : PG_17 port map( p1 => psignal_0_23_port, g1 => 
                           gsignal_0_23_port, p2 => psignal_0_22_port, g2 => 
                           gsignal_0_22_port, p_Out => psignal_1_23_port, g_Out
                           => gsignal_1_23_port);
   PGelements_0_25 : PG_16 port map( p1 => psignal_0_25_port, g1 => 
                           gsignal_0_25_port, p2 => psignal_0_24_port, g2 => 
                           gsignal_0_24_port, p_Out => psignal_1_25_port, g_Out
                           => gsignal_1_25_port);
   PGelements_0_27 : PG_15 port map( p1 => psignal_0_27_port, g1 => 
                           gsignal_0_27_port, p2 => psignal_0_26_port, g2 => 
                           gsignal_0_26_port, p_Out => psignal_1_27_port, g_Out
                           => gsignal_1_27_port);
   PGelements_0_29 : PG_14 port map( p1 => psignal_0_29_port, g1 => 
                           gsignal_0_29_port, p2 => psignal_0_28_port, g2 => 
                           gsignal_0_28_port, p_Out => psignal_1_29_port, g_Out
                           => gsignal_1_29_port);
   PGelements_0_31 : PG_13 port map( p1 => psignal_0_31_port, g1 => 
                           gsignal_0_31_port, p2 => psignal_0_30_port, g2 => 
                           gsignal_0_30_port, p_Out => psignal_1_31_port, g_Out
                           => gsignal_1_31_port);
   g0_1_3 : G_8 port map( p1 => psignal_1_3_port, g1 => gsignal_1_3_port, g2 =>
                           gsignal_1_1_port, g_Out => n7);
   PGelements_1_7 : PG_12 port map( p1 => psignal_1_7_port, g1 => 
                           gsignal_1_7_port, p2 => psignal_1_5_port, g2 => 
                           gsignal_1_5_port, p_Out => psignal_2_7_port, g_Out 
                           => gsignal_2_7_port);
   PGelements_1_11 : PG_11 port map( p1 => psignal_1_11_port, g1 => 
                           gsignal_1_11_port, p2 => psignal_1_9_port, g2 => 
                           gsignal_1_9_port, p_Out => psignal_2_11_port, g_Out 
                           => gsignal_2_11_port);
   PGelements_1_15 : PG_10 port map( p1 => psignal_1_15_port, g1 => 
                           gsignal_1_15_port, p2 => psignal_1_13_port, g2 => 
                           gsignal_1_13_port, p_Out => psignal_2_15_port, g_Out
                           => gsignal_2_15_port);
   PGelements_1_19 : PG_9 port map( p1 => psignal_1_19_port, g1 => 
                           gsignal_1_19_port, p2 => psignal_1_17_port, g2 => 
                           gsignal_1_17_port, p_Out => psignal_2_19_port, g_Out
                           => gsignal_2_19_port);
   PGelements_1_23 : PG_8 port map( p1 => psignal_1_23_port, g1 => 
                           gsignal_1_23_port, p2 => psignal_1_21_port, g2 => 
                           gsignal_1_21_port, p_Out => psignal_2_23_port, g_Out
                           => gsignal_2_23_port);
   PGelements_1_27 : PG_7 port map( p1 => psignal_1_27_port, g1 => 
                           gsignal_1_27_port, p2 => psignal_1_25_port, g2 => 
                           gsignal_1_25_port, p_Out => psignal_2_27_port, g_Out
                           => gsignal_2_27_port);
   PGelements_1_31 : PG_6 port map( p1 => psignal_1_31_port, g1 => 
                           gsignal_1_31_port, p2 => psignal_1_29_port, g2 => 
                           gsignal_1_29_port, p_Out => psignal_2_31_port, g_Out
                           => gsignal_2_31_port);
   g0_2_7 : G_7 port map( p1 => psignal_2_7_port, g1 => gsignal_2_7_port, g2 =>
                           n7, g_Out => n6);
   PGelements_2_15 : PG_5 port map( p1 => psignal_2_15_port, g1 => 
                           gsignal_2_15_port, p2 => psignal_2_11_port, g2 => 
                           gsignal_2_11_port, p_Out => psignal_3_15_port, g_Out
                           => gsignal_3_15_port);
   PGelements_2_23 : PG_4 port map( p1 => psignal_2_23_port, g1 => 
                           gsignal_2_23_port, p2 => psignal_2_19_port, g2 => 
                           gsignal_2_19_port, p_Out => psignal_3_23_port, g_Out
                           => gsignal_3_23_port);
   PGelements_2_31 : PG_3 port map( p1 => psignal_2_31_port, g1 => 
                           gsignal_2_31_port, p2 => psignal_2_27_port, g2 => 
                           gsignal_2_27_port, p_Out => psignal_3_31_port, g_Out
                           => gsignal_3_31_port);
   g1_3_11 : G_6 port map( p1 => psignal_2_11_port, g1 => gsignal_2_11_port, g2
                           => cout_1_port, g_Out => cout_2_port);
   g1_3_15 : G_5 port map( p1 => psignal_3_15_port, g1 => gsignal_3_15_port, g2
                           => n6, g_Out => n3);
   pg1_3_27 : PG_2 port map( p1 => psignal_2_27_port, g1 => gsignal_2_27_port, 
                           p2 => psignal_3_15_port, g2 => gsignal_3_15_port, 
                           p_Out => psignal_4_27_port, g_Out => 
                           gsignal_4_27_port);
   pg1_3_31 : PG_1 port map( p1 => psignal_3_31_port, g1 => gsignal_3_31_port, 
                           p2 => psignal_3_15_port, g2 => gsignal_3_15_port, 
                           p_Out => psignal_4_31_port, g_Out => 
                           gsignal_4_31_port);
   g1_4_19 : G_4 port map( p1 => psignal_2_19_port, g1 => gsignal_2_19_port, g2
                           => n3, g_Out => cout_4_port);
   g1_4_23 : G_3 port map( p1 => psignal_3_23_port, g1 => gsignal_3_23_port, g2
                           => n3, g_Out => cout_5_port);
   g1_4_27 : G_2 port map( p1 => psignal_4_27_port, g1 => gsignal_4_27_port, g2
                           => n3, g_Out => cout_6_port);
   g1_4_31 : G_1 port map( p1 => psignal_4_31_port, g1 => gsignal_4_31_port, g2
                           => n3, g_Out => cout_7_port);
   U1 : BUF_X1 port map( A => n7, Z => cout_0_port);
   U3 : BUF_X2 port map( A => n6, Z => cout_1_port);
   U4 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => g0);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity SHIFTER_M32_N5_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (31 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_M32_N5_DW_rash_0;

architecture SYN_mx2 of SHIFTER_M32_N5_DW_rash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X4
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n201, n202, n203, n204, n205, n206, n208, n209, n210, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n240, n241, n242, n243, n244, n245, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n260, n261, n263, n265, 
      n266, n268, n272, n273, n279, n280, n283, n286, n287, n290, n291, n294, 
      n295, n298, n299, n302, n303, n305, n306, n309, n310, n314, n315, n316, 
      n317, n318, n321, n322, n325, n326, n327, n329, n330, n331, n332, n334, 
      n335, n336, n337, n338, n341, n342, n343, n344, n347, n348, n350, n351, 
      n352, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n371, n372, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n385, n387, n388, n424, n477, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n566, 
      n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698 : 
      std_logic;

begin
   
   U93 : NAND3_X1 port map( A1 => n585, A2 => n696, A3 => n102, ZN => n100);
   U96 : MUX2_X1 port map( A => n109, B => n110, S => n111, Z => n108);
   U98 : MUX2_X1 port map( A => n115, B => n116, S => n111, Z => n114);
   U100 : MUX2_X1 port map( A => n119, B => n120, S => n111, Z => n118);
   U102 : MUX2_X1 port map( A => n123, B => n124, S => n111, Z => n122);
   U104 : MUX2_X1 port map( A => n127, B => n128, S => n111, Z => n126);
   U106 : MUX2_X1 port map( A => n577, B => n131, S => n111, Z => n129);
   U109 : NAND3_X1 port map( A1 => n136, A2 => n137, A3 => n132, ZN => n135);
   U132 : NAND3_X1 port map( A1 => n585, A2 => n696, A3 => n170, ZN => n177);
   U141 : MUX2_X1 port map( A => n182, B => n183, S => n111, Z => n181);
   U197 : NAND3_X1 port map( A1 => n136, A2 => n137, A3 => n206, ZN => n208);
   U244 : MUX2_X1 port map( A => n189, B => n190, S => n111, Z => n227);
   U23 : NAND3_X1 port map( A1 => n290, A2 => n291, A3 => n204, ZN => n263);
   U46 : NAND3_X1 port map( A1 => n351, A2 => n350, A3 => n197, ZN => n142);
   U59 : NAND3_X1 port map( A1 => n279, A2 => n280, A3 => n212, ZN => n162);
   U71 : NAND3_X1 port map( A1 => n286, A2 => n287, A3 => n198, ZN => n144);
   U76 : NAND3_X1 port map( A1 => n290, A2 => n291, A3 => n204, ZN => n149);
   U81 : NAND3_X1 port map( A1 => n294, A2 => n295, A3 => n233, ZN => n152);
   U86 : NAND3_X1 port map( A1 => n298, A2 => n299, A3 => n225, ZN => n176);
   U94 : NAND3_X1 port map( A1 => n302, A2 => n303, A3 => n236, ZN => n158);
   U107 : NAND3_X1 port map( A1 => n305, A2 => n306, A3 => n199, ZN => n148);
   U122 : NAND3_X1 port map( A1 => n314, A2 => n315, A3 => n232, ZN => n157);
   U130 : NAND3_X1 port map( A1 => n224, A2 => n338, A3 => n337, ZN => n321);
   U138 : NAND3_X1 port map( A1 => n325, A2 => n326, A3 => n203, ZN => n145);
   U154 : NAND3_X1 port map( A1 => n337, A2 => n338, A3 => n224, ZN => n172);
   U170 : NAND3_X1 port map( A1 => n347, A2 => n348, A3 => n223, ZN => n169);
   U182 : NAND3_X1 port map( A1 => n358, A2 => n359, A3 => n217, ZN => n164);
   U190 : NAND3_X1 port map( A1 => n365, A2 => n366, A3 => n216, ZN => n167);
   U193 : NAND3_X1 port map( A1 => n367, A2 => n368, A3 => n235, ZN => n150);
   U200 : NAND3_X1 port map( A1 => n371, A2 => n372, A3 => n202, ZN => n141);
   U208 : NAND3_X1 port map( A1 => n215, A2 => n380, A3 => n379, ZN => n163);
   U373 : NAND3_X1 port map( A1 => SH(15), A2 => SH(14), A3 => SH(16), ZN => 
                           n506);
   U281 : NAND2_X2 port map( A1 => SH(4), A2 => n228, ZN => n111);
   U3 : BUF_X1 port map( A => n273, Z => n596);
   U4 : CLKBUF_X1 port map( A => n240, Z => n566);
   U5 : CLKBUF_X3 port map( A => n272, Z => n639);
   U6 : CLKBUF_X2 port map( A => n272, Z => n638);
   U7 : OAI221_X1 port map( B1 => n616, B2 => n680, C1 => n620, C2 => n676, A 
                           => n219, ZN => n175);
   U8 : BUF_X2 port map( A => n261, Z => n641);
   U9 : OR2_X1 port map( A1 => n694, A2 => n218, ZN => n113);
   U10 : NOR3_X1 port map( A1 => n588, A2 => n589, A3 => n590, ZN => n131);
   U11 : AND2_X1 port map( A1 => n164, A2 => n643, ZN => n330);
   U12 : AND3_X1 port map( A1 => n481, A2 => n482, A3 => n180, ZN => n105);
   U13 : AOI22_X1 port map( A1 => A(30), A2 => n637, B1 => n639, B2 => A(31), 
                           ZN => n117);
   U14 : BUF_X2 port map( A => n261, Z => n643);
   U15 : NOR3_X1 port map( A1 => n608, A2 => n609, A3 => n655, ZN => n134);
   U16 : CLKBUF_X1 port map( A => n240, Z => n567);
   U17 : AND2_X2 port map( A1 => n344, A2 => SH(1), ZN => n383);
   U18 : BUF_X1 port map( A => n155, Z => n568);
   U19 : CLKBUF_X1 port map( A => n145, Z => n569);
   U20 : AND4_X1 port map( A1 => n247, A2 => SH(22), A3 => SH(20), A4 => SH(21)
                           , ZN => n244);
   U21 : OR2_X1 port map( A1 => n268, A2 => n690, ZN => n570);
   U22 : NAND3_X1 port map( A1 => n317, A2 => n318, A3 => n221, ZN => n571);
   U24 : OAI221_X1 port map( B1 => n594, B2 => n689, C1 => n619, C2 => n684, A 
                           => n231, ZN => n572);
   U25 : AOI22_X1 port map( A1 => A(24), A2 => n638, B1 => A(25), B2 => n631, 
                           ZN => n573);
   U26 : BUF_X1 port map( A => n273, Z => n595);
   U27 : NAND2_X1 port map( A1 => n155, A2 => n627, ZN => n574);
   U28 : NAND2_X1 port map( A1 => n158, A2 => n641, ZN => n575);
   U29 : NAND2_X1 port map( A1 => n574, A2 => n575, ZN => n576);
   U30 : NOR2_X1 port map( A1 => n424, A2 => n576, ZN => n577);
   U31 : BUF_X2 port map( A => n385, Z => n578);
   U32 : NAND2_X1 port map( A1 => n624, A2 => A(15), ZN => n336);
   U33 : AOI222_X4 port map( A1 => n578, A2 => A(1), B1 => n638, B2 => A(0), C1
                           => n598, C2 => A(2), ZN => n106);
   U34 : MUX2_X1 port map( A => n160, B => n159, S => n196, Z => n136);
   U35 : OAI221_X1 port map( B1 => n693, B2 => n94, C1 => n691, C2 => n93, A =>
                           n570, ZN => B(7));
   U36 : AND3_X1 port map( A1 => n336, A2 => n335, A3 => n230, ZN => n266);
   U37 : OAI22_X1 port map( A1 => n615, A2 => n579, B1 => n106, B2 => n580, ZN 
                           => n581);
   U38 : INV_X1 port map( A => n600, ZN => n579);
   U39 : INV_X1 port map( A => n261, ZN => n580);
   U40 : INV_X1 port map( A => n581, ZN => n94);
   U41 : NAND2_X1 port map( A1 => n584, A2 => n566, ZN => n273);
   U42 : OAI22_X1 port map( A1 => n266, A2 => n615, B1 => n582, B2 => n614, ZN 
                           => n668);
   U43 : INV_X1 port map( A => n153, ZN => n582);
   U44 : NAND3_X1 port map( A1 => n336, A2 => n335, A3 => n230, ZN => n154);
   U45 : NAND3_X1 port map( A1 => n209, A2 => n343, A3 => n342, ZN => n159);
   U47 : NAND3_X1 port map( A1 => n364, A2 => n363, A3 => n362, ZN => n648);
   U48 : BUF_X1 port map( A => n161, Z => n583);
   U49 : AND2_X1 port map( A1 => n165, A2 => n612, ZN => n268);
   U50 : INV_X1 port map( A => n383, ZN => n584);
   U51 : CLKBUF_X1 port map( A => n101, Z => n585);
   U52 : NAND3_X1 port map( A1 => n331, A2 => n332, A3 => n210, ZN => n586);
   U53 : NAND3_X1 port map( A1 => n294, A2 => n295, A3 => n233, ZN => n587);
   U54 : AND2_X1 port map( A1 => n152, A2 => n642, ZN => n588);
   U55 : AND2_X1 port map( A1 => n153, A2 => n626, ZN => n589);
   U56 : AND2_X1 port map( A1 => n157, A2 => n628, ZN => n590);
   U57 : OR2_X1 port map( A1 => n567, A2 => n698, ZN => n591);
   U58 : OR2_X1 port map( A1 => n567, A2 => n698, ZN => n334);
   U60 : NAND3_X1 port map( A1 => n358, A2 => n359, A3 => n217, ZN => n592);
   U61 : BUF_X1 port map( A => n240, Z => n604);
   U62 : CLKBUF_X1 port map( A => SH(17), Z => n593);
   U63 : INV_X1 port map( A => n165, ZN => n660);
   U64 : CLKBUF_X1 port map( A => n273, Z => n594);
   U65 : CLKBUF_X3 port map( A => n272, Z => n640);
   U66 : INV_X1 port map( A => n334, ZN => n597);
   U67 : INV_X1 port map( A => n591, ZN => n598);
   U68 : INV_X1 port map( A => n591, ZN => n599);
   U69 : INV_X1 port map( A => n334, ZN => n624);
   U70 : NAND3_X1 port map( A1 => n279, A2 => n280, A3 => n212, ZN => n600);
   U72 : OAI221_X1 port map( B1 => n616, B2 => n659, C1 => n656, C2 => n620, A 
                           => n214, ZN => n601);
   U73 : NAND3_X1 port map( A1 => n215, A2 => n380, A3 => n379, ZN => n602);
   U74 : CLKBUF_X1 port map( A => n142, Z => n603);
   U75 : AND2_X1 port map( A1 => n148, A2 => n628, ZN => n605);
   U77 : AND2_X1 port map( A1 => n144, A2 => n642, ZN => n606);
   U78 : AND2_X1 port map( A1 => n137, A2 => n101, ZN => n607);
   U79 : NOR3_X1 port map( A1 => n605, A2 => n606, A3 => n607, ZN => n128);
   U80 : BUF_X1 port map( A => n385, Z => n630);
   U82 : AND2_X1 port map( A1 => n592, A2 => n627, ZN => n608);
   U83 : AND2_X1 port map( A1 => n167, A2 => n641, ZN => n609);
   U84 : AND2_X1 port map( A1 => n240, A2 => n383, ZN => n385);
   U85 : AND4_X1 port map( A1 => n249, A2 => SH(9), A3 => SH(7), A4 => SH(8), 
                           ZN => n610);
   U87 : CLKBUF_X1 port map( A => SH(28), Z => n611);
   U88 : AND4_X1 port map( A1 => n249, A2 => SH(9), A3 => SH(7), A4 => SH(8), 
                           ZN => n242);
   U89 : MUX2_X2 port map( A => n142, B => n143, S => n196, Z => n101);
   U90 : NOR2_X1 port map( A1 => n330, A2 => n329, ZN => n612);
   U91 : BUF_X2 port map( A => n385, Z => n613);
   U92 : INV_X4 port map( A => n102, ZN => n693);
   U95 : INV_X2 port map( A => n132, ZN => n690);
   U97 : INV_X2 port map( A => n614, ZN => n634);
   U99 : INV_X1 port map( A => n614, ZN => n633);
   U101 : INV_X1 port map( A => n170, ZN => n692);
   U103 : NAND2_X1 port map( A1 => n170, A2 => n628, ZN => n179);
   U105 : NAND2_X1 port map( A1 => n132, A2 => n633, ZN => n112);
   U108 : INV_X1 port map( A => n615, ZN => n628);
   U110 : OAI222_X1 port map( A1 => n89, A2 => n693, B1 => n91, B2 => n692, C1 
                           => n90, C2 => n690, ZN => B(24));
   U111 : NOR2_X1 port map( A1 => n107, A2 => n695, ZN => n132);
   U112 : INV_X1 port map( A => n206, ZN => n691);
   U113 : BUF_X2 port map( A => n387, Z => n625);
   U114 : NOR2_X1 port map( A1 => n113, A2 => n695, ZN => n170);
   U115 : BUF_X2 port map( A => n385, Z => n631);
   U116 : BUF_X2 port map( A => n387, Z => n626);
   U117 : OAI222_X1 port map( A1 => n103, A2 => n691, B1 => n683, B2 => n104, 
                           C1 => n105, C2 => n690, ZN => B(4));
   U118 : OAI222_X1 port map( A1 => n86, A2 => n690, B1 => n87, B2 => n691, C1 
                           => n88, C2 => n693, ZN => B(9));
   U119 : OAI221_X1 port map( B1 => n98, B2 => n691, C1 => n99, C2 => n690, A 
                           => n100, ZN => B(5));
   U120 : OAI222_X1 port map( A1 => n577, A2 => n690, B1 => n644, B2 => n191, 
                           C1 => n131, C2 => n693, ZN => B(12));
   U121 : OAI222_X1 port map( A1 => n138, A2 => n690, B1 => n140, B2 => n691, 
                           C1 => n139, C2 => n693, ZN => B(10));
   U123 : BUF_X2 port map( A => n261, Z => n642);
   U124 : BUF_X2 port map( A => n387, Z => n627);
   U125 : BUF_X2 port map( A => n385, Z => n632);
   U126 : OR2_X2 port map( A1 => n697, A2 => n696, ZN => n614);
   U127 : NAND2_X1 port map( A1 => n102, A2 => n628, ZN => n104);
   U128 : NOR3_X1 port map( A1 => n381, A2 => n382, A3 => n651, ZN => n119);
   U129 : NAND2_X1 port map( A1 => n206, A2 => n633, ZN => n191);
   U131 : OAI222_X1 port map( A1 => n92, A2 => n693, B1 => n94, B2 => n692, C1 
                           => n93, C2 => n690, ZN => B(23));
   U133 : OAI222_X1 port map( A1 => n86, A2 => n693, B1 => n88, B2 => n692, C1 
                           => n87, C2 => n690, ZN => B(25));
   U134 : INV_X1 port map( A => n143, ZN => n688);
   U135 : OAI222_X1 port map( A1 => n95, A2 => n690, B1 => n96, B2 => n691, C1 
                           => n97, C2 => n693, ZN => B(6));
   U136 : OAI222_X1 port map( A1 => n183, A2 => n693, B1 => n688, B2 => n179, 
                           C1 => n182, C2 => n690, ZN => B(17));
   U137 : OAI222_X1 port map( A1 => n138, A2 => n693, B1 => n139, B2 => n692, 
                           C1 => n140, C2 => n690, ZN => B(26));
   U139 : OAI221_X1 port map( B1 => n99, B2 => n693, C1 => n98, C2 => n690, A 
                           => n177, ZN => B(21));
   U140 : AND3_X1 port map( A1 => n192, A2 => n674, A3 => n679, ZN => n352);
   U142 : INV_X1 port map( A => n377, ZN => n679);
   U143 : INV_X1 port map( A => n378, ZN => n674);
   U144 : INV_X1 port map( A => n160, ZN => n645);
   U145 : NOR2_X1 port map( A1 => n107, A2 => n227, ZN => B(0));
   U146 : AOI222_X1 port map( A1 => n647, A2 => n643, B1 => n571, B2 => n626, 
                           C1 => n169, C2 => n633, ZN => n96);
   U147 : AOI222_X1 port map( A1 => n171, A2 => n643, B1 => n687, B2 => n626, 
                           C1 => n175, C2 => n628, ZN => n139);
   U148 : AOI222_X1 port map( A1 => n159, A2 => n626, B1 => n643, B2 => n160, 
                           C1 => n161, C2 => n633, ZN => n93);
   U149 : AOI222_X1 port map( A1 => n151, A2 => n642, B1 => n150, B2 => n626, 
                           C1 => n158, C2 => n633, ZN => n103);
   U150 : AOI222_X1 port map( A1 => n648, A2 => n642, B1 => n141, B2 => n626, 
                           C1 => n263, C2 => n633, ZN => n98);
   U151 : OAI22_X1 port map( A1 => n615, A2 => n265, B1 => n614, B2 => n266, ZN
                           => n424);
   U152 : AND3_X1 port map( A1 => n367, A2 => n368, A3 => n235, ZN => n265);
   U153 : AOI221_X1 port map( B1 => n152, B2 => n627, C1 => n157, C2 => n641, A
                           => n668, ZN => n190);
   U155 : NOR2_X1 port map( A1 => n113, A2 => n111, ZN => n102);
   U156 : AOI22_X1 port map( A1 => n571, A2 => n633, B1 => n647, B2 => n626, ZN
                           => n140);
   U157 : AOI22_X1 port map( A1 => n141, A2 => n633, B1 => n648, B2 => n626, ZN
                           => n87);
   U158 : AOI22_X1 port map( A1 => n150, A2 => n633, B1 => n151, B2 => n626, ZN
                           => n90);
   U159 : AOI22_X1 port map( A1 => n171, A2 => n628, B1 => n687, B2 => n642, ZN
                           => n97);
   U160 : NOR2_X1 port map( A1 => n107, A2 => n111, ZN => n206);
   U161 : NAND2_X1 port map( A1 => n218, A2 => n694, ZN => n107);
   U162 : NOR2_X1 port map( A1 => n635, A2 => n646, ZN => n160);
   U163 : AOI22_X1 port map( A1 => n634, A2 => n686, B1 => n629, B2 => n602, ZN
                           => n192);
   U164 : OAI222_X1 port map( A1 => n89, A2 => n690, B1 => n90, B2 => n691, C1 
                           => n91, C2 => n693, ZN => B(8));
   U165 : OAI22_X1 port map( A1 => n125, A2 => n112, B1 => n126, B2 => n113, ZN
                           => B(29));
   U166 : INV_X1 port map( A => n193, ZN => n649);
   U167 : AOI22_X1 port map( A1 => n634, A2 => n592, B1 => n629, B2 => n159, ZN
                           => n193);
   U168 : NOR2_X1 port map( A1 => n689, A2 => n621, ZN => n143);
   U169 : INV_X1 port map( A => n106, ZN => n686);
   U171 : AND3_X1 port map( A1 => n483, A2 => n484, A3 => n178, ZN => n99);
   U172 : NAND2_X1 port map( A1 => n569, A2 => n642, ZN => n484);
   U173 : NAND2_X1 port map( A1 => n148, A2 => n625, ZN => n483);
   U174 : AOI22_X1 port map( A1 => n634, A2 => n144, B1 => n628, B2 => n146, ZN
                           => n178);
   U175 : AOI22_X1 port map( A1 => n634, A2 => n602, B1 => n601, B2 => n628, ZN
                           => n213);
   U176 : AND3_X1 port map( A1 => n495, A2 => n496, A3 => n201, ZN => n127);
   U177 : NAND2_X1 port map( A1 => n149, A2 => n641, ZN => n496);
   U178 : NAND2_X1 port map( A1 => n146, A2 => n625, ZN => n495);
   U179 : AOI22_X1 port map( A1 => n634, A2 => n145, B1 => n629, B2 => n141, ZN
                           => n201);
   U180 : NAND2_X1 port map( A1 => n157, A2 => n625, ZN => n481);
   U181 : AOI22_X1 port map( A1 => n634, A2 => n587, B1 => n155, B2 => n628, ZN
                           => n180);
   U183 : AND3_X1 port map( A1 => n186, A2 => n260, A3 => n477, ZN => n124);
   U184 : NAND2_X1 port map( A1 => n172, A2 => n642, ZN => n260);
   U185 : NAND2_X1 port map( A1 => n175, A2 => n625, ZN => n477);
   U186 : AOI22_X1 port map( A1 => n634, A2 => n171, B1 => n629, B2 => n173, ZN
                           => n186);
   U187 : AND3_X1 port map( A1 => n487, A2 => n488, A3 => n174, ZN => n95);
   U188 : NAND2_X1 port map( A1 => n173, A2 => n641, ZN => n488);
   U189 : NAND2_X1 port map( A1 => n321, A2 => n625, ZN => n487);
   U191 : AOI22_X1 port map( A1 => n175, A2 => n633, B1 => n628, B2 => n176, ZN
                           => n174);
   U192 : OAI22_X1 port map( A1 => n108, A2 => n107, B1 => n104, B2 => n106, ZN
                           => B(3));
   U194 : OR2_X1 port map( A1 => n196, A2 => n137, ZN => n615);
   U195 : NOR3_X1 port map( A1 => n376, A2 => n375, A3 => n374, ZN => n109);
   U196 : AND2_X1 port map( A1 => n192, A2 => n310, ZN => n116);
   U198 : NOR3_X1 port map( A1 => n356, A2 => n357, A3 => n649, ZN => n115);
   U199 : NOR2_X1 port map( A1 => n378, A2 => n377, ZN => n310);
   U201 : INV_X1 port map( A => n121, ZN => n687);
   U202 : INV_X1 port map( A => n117, ZN => n647);
   U203 : INV_X1 port map( A => n151, ZN => n644);
   U204 : INV_X1 port map( A => n111, ZN => n695);
   U205 : AND3_X1 port map( A1 => n485, A2 => n486, A3 => n147, ZN => n86);
   U206 : NAND2_X1 port map( A1 => n569, A2 => n625, ZN => n485);
   U207 : NAND2_X1 port map( A1 => n146, A2 => n642, ZN => n486);
   U209 : AOI22_X1 port map( A1 => n634, A2 => n148, B1 => n629, B2 => n149, ZN
                           => n147);
   U210 : AND3_X1 port map( A1 => n489, A2 => n490, A3 => n156, ZN => n89);
   U211 : NAND2_X1 port map( A1 => n568, A2 => n641, ZN => n490);
   U212 : AOI22_X1 port map( A1 => n634, A2 => n157, B1 => n628, B2 => n158, ZN
                           => n156);
   U213 : AND3_X1 port map( A1 => n491, A2 => n492, A3 => n222, ZN => n138);
   U214 : NAND2_X1 port map( A1 => n173, A2 => n625, ZN => n491);
   U215 : NAND2_X1 port map( A1 => n176, A2 => n641, ZN => n492);
   U216 : AOI22_X1 port map( A1 => n634, A2 => n321, B1 => n629, B2 => n169, ZN
                           => n222);
   U217 : AND2_X1 port map( A1 => n601, A2 => n627, ZN => n375);
   U218 : AND2_X1 port map( A1 => n169, A2 => n643, ZN => n382);
   U219 : AND2_X1 port map( A1 => n176, A2 => n627, ZN => n381);
   U220 : OAI222_X1 port map( A1 => n95, A2 => n693, B1 => n97, B2 => n692, C1 
                           => n96, C2 => n690, ZN => B(22));
   U221 : OAI22_X1 port map( A1 => n121, A2 => n104, B1 => n107, B2 => n122, ZN
                           => B(2));
   U222 : OAI22_X1 port map( A1 => n644, A2 => n112, B1 => n113, B2 => n129, ZN
                           => B(28));
   U223 : AND2_X1 port map( A1 => n162, A2 => n627, ZN => n377);
   U224 : AND2_X1 port map( A1 => n166, A2 => n643, ZN => n378);
   U225 : INV_X1 port map( A => n195, ZN => n651);
   U226 : AND3_X1 port map( A1 => n493, A2 => n494, A3 => n185, ZN => n123);
   U227 : NAND2_X1 port map( A1 => n168, A2 => n641, ZN => n494);
   U228 : NAND2_X1 port map( A1 => n169, A2 => n625, ZN => n493);
   U229 : AOI22_X1 port map( A1 => n634, A2 => n176, B1 => n629, B2 => n647, ZN
                           => n185);
   U230 : AND3_X1 port map( A1 => n497, A2 => n498, A3 => n188, ZN => n183);
   U231 : NAND2_X1 port map( A1 => n144, A2 => n625, ZN => n497);
   U232 : NAND2_X1 port map( A1 => n148, A2 => n641, ZN => n498);
   U233 : AND3_X1 port map( A1 => n499, A2 => n500, A3 => n184, ZN => n110);
   U234 : NAND2_X1 port map( A1 => n586, A2 => n625, ZN => n499);
   U235 : NAND2_X1 port map( A1 => n602, A2 => n641, ZN => n500);
   U236 : AND3_X1 port map( A1 => n503, A2 => n504, A3 => n194, ZN => n120);
   U237 : NAND2_X1 port map( A1 => n171, A2 => n625, ZN => n503);
   U238 : NAND2_X1 port map( A1 => n175, A2 => n641, ZN => n504);
   U239 : AOI22_X1 port map( A1 => n634, A2 => n687, B1 => n629, B2 => n172, ZN
                           => n194);
   U240 : AND2_X1 port map( A1 => n583, A2 => n643, ZN => n357);
   U241 : AND2_X1 port map( A1 => n327, A2 => n187, ZN => n182);
   U242 : AOI22_X1 port map( A1 => n634, A2 => n146, B1 => n629, B2 => n648, ZN
                           => n187);
   U243 : NOR2_X1 port map( A1 => n360, A2 => n361, ZN => n327);
   U245 : AND2_X1 port map( A1 => n263, A2 => n627, ZN => n360);
   U246 : AND3_X1 port map( A1 => n501, A2 => n502, A3 => n234, ZN => n189);
   U247 : NAND2_X1 port map( A1 => n151, A2 => n628, ZN => n502);
   U248 : NAND2_X1 port map( A1 => n568, A2 => n633, ZN => n501);
   U249 : AOI22_X1 port map( A1 => n626, A2 => n158, B1 => n643, B2 => n150, ZN
                           => n234);
   U250 : AND2_X1 port map( A1 => n163, A2 => n627, ZN => n329);
   U251 : OAI222_X1 port map( A1 => n316, A2 => n690, B1 => n117, B2 => n191, 
                           C1 => n693, C2 => n120, ZN => B(14));
   U252 : NOR3_X1 port map( A1 => n381, A2 => n382, A3 => n651, ZN => n316);
   U253 : OAI222_X1 port map( A1 => n105, A2 => n693, B1 => n683, B2 => n179, 
                           C1 => n103, C2 => n690, ZN => B(20));
   U254 : OAI222_X1 port map( A1 => n124, A2 => n693, B1 => n121, B2 => n179, 
                           C1 => n123, C2 => n690, ZN => B(18));
   U255 : INV_X1 port map( A => n196, ZN => n697);
   U256 : AND2_X1 port map( A1 => n141, A2 => n643, ZN => n361);
   U257 : OAI222_X1 port map( A1 => n110, A2 => n693, B1 => n106, B2 => n179, 
                           C1 => n341, C2 => n690, ZN => B(19));
   U258 : NOR3_X1 port map( A1 => n376, A2 => n375, A3 => n374, ZN => n341);
   U259 : OR2_X1 port map( A1 => n654, A2 => n620, ZN => n368);
   U260 : OR2_X1 port map( A1 => n623, A2 => n671, ZN => n338);
   U261 : OR2_X1 port map( A1 => n622, A2 => n658, ZN => n291);
   U262 : OR2_X1 port map( A1 => n635, A2 => n675, ZN => n337);
   U263 : OAI221_X1 port map( B1 => n616, B2 => n685, C1 => n618, C2 => n681, A
                           => n220, ZN => n171);
   U264 : OAI221_X1 port map( B1 => n635, B2 => n666, C1 => n619, C2 => n663, A
                           => n205, ZN => n146);
   U265 : AOI22_X1 port map( A1 => A(18), A2 => n640, B1 => A(19), B2 => n578, 
                           ZN => n205);
   U266 : OAI221_X1 port map( B1 => n616, B2 => n667, C1 => n620, C2 => n664, A
                           => n238, ZN => n155);
   U267 : AOI22_X1 port map( A1 => A(17), A2 => n640, B1 => A(18), B2 => n631, 
                           ZN => n238);
   U268 : AOI22_X1 port map( A1 => A(7), A2 => n639, B1 => A(8), B2 => n632, ZN
                           => n219);
   U269 : OAI221_X1 port map( B1 => n594, B2 => n653, C1 => n646, C2 => n622, A
                           => n237, ZN => n151);
   U270 : AOI22_X1 port map( A1 => A(29), A2 => n639, B1 => n630, B2 => A(30), 
                           ZN => n237);
   U271 : OR2_X1 port map( A1 => n622, A2 => n672, ZN => n306);
   U272 : AOI22_X1 port map( A1 => A(21), A2 => n640, B1 => A(22), B2 => n632, 
                           ZN => n236);
   U273 : OR2_X1 port map( A1 => n618, A2 => n659, ZN => n303);
   U274 : AOI22_X1 port map( A1 => A(6), A2 => n640, B1 => A(7), B2 => n578, ZN
                           => n198);
   U275 : OR2_X1 port map( A1 => n619, A2 => n677, ZN => n287);
   U276 : AOI22_X1 port map( A1 => A(12), A2 => n638, B1 => A(13), B2 => n578, 
                           ZN => n215);
   U277 : OR2_X1 port map( A1 => n621, A2 => n670, ZN => n380);
   U278 : OR2_X1 port map( A1 => n596, A2 => n665, ZN => n298);
   U279 : AOI22_X1 port map( A1 => A(19), A2 => n640, B1 => A(20), B2 => n631, 
                           ZN => n225);
   U280 : OR2_X1 port map( A1 => n619, A2 => n662, ZN => n299);
   U282 : AOI22_X1 port map( A1 => A(26), A2 => n639, B1 => A(27), B2 => n631, 
                           ZN => n202);
   U283 : OR2_X1 port map( A1 => n623, A2 => n653, ZN => n372);
   U284 : OR2_X1 port map( A1 => n622, A2 => n673, ZN => n315);
   U285 : OR2_X1 port map( A1 => n616, A2 => n671, ZN => n325);
   U286 : AOI22_X1 port map( A1 => A(14), A2 => n639, B1 => A(15), B2 => n631, 
                           ZN => n203);
   U287 : OR2_X1 port map( A1 => n619, A2 => n667, ZN => n326);
   U288 : AOI22_X1 port map( A1 => A(23), A2 => n640, B1 => A(24), B2 => n578, 
                           ZN => n223);
   U289 : OR2_X1 port map( A1 => n635, A2 => n661, ZN => n347);
   U290 : OR2_X1 port map( A1 => n657, A2 => n620, ZN => n348);
   U291 : AOI22_X1 port map( A1 => A(5), A2 => n640, B1 => A(6), B2 => n578, ZN
                           => n233);
   U292 : OR2_X1 port map( A1 => n619, A2 => n678, ZN => n295);
   U293 : AOI22_X1 port map( A1 => A(16), A2 => n638, B1 => n632, B2 => A(17), 
                           ZN => n217);
   U294 : OR2_X1 port map( A1 => n618, A2 => n665, ZN => n359);
   U295 : AOI22_X1 port map( A1 => A(20), A2 => n638, B1 => A(21), B2 => n613, 
                           ZN => n216);
   U296 : OR2_X1 port map( A1 => n622, A2 => n661, ZN => n366);
   U297 : AOI22_X1 port map( A1 => A(28), A2 => n638, B1 => A(29), B2 => n613, 
                           ZN => n209);
   U298 : OR2_X1 port map( A1 => n650, A2 => n617, ZN => n343);
   U299 : OR2_X1 port map( A1 => n623, A2 => n680, ZN => n280);
   U300 : AOI22_X1 port map( A1 => n640, A2 => A(25), B1 => A(26), B2 => n630, 
                           ZN => n235);
   U301 : AOI21_X1 port map( B1 => n250, B2 => n694, A => SH(5), ZN => n218);
   U302 : NAND4_X1 port map( A1 => n251, A2 => n252, A3 => n253, A4 => n254, ZN
                           => n250);
   U303 : AOI22_X1 port map( A1 => A(13), A2 => n639, B1 => A(14), B2 => n578, 
                           ZN => n230);
   U304 : AOI22_X1 port map( A1 => A(22), A2 => n639, B1 => A(23), B2 => n630, 
                           ZN => n204);
   U305 : OAI221_X1 port map( B1 => n616, B2 => n659, C1 => n656, C2 => n620, A
                           => n573, ZN => n161);
   U306 : AOI22_X1 port map( A1 => A(24), A2 => n638, B1 => A(25), B2 => n631, 
                           ZN => n214);
   U307 : AOI22_X1 port map( A1 => A(11), A2 => n640, B1 => A(12), B2 => n630, 
                           ZN => n224);
   U308 : NAND2_X1 port map( A1 => SH(3), A2 => n228, ZN => n137);
   U309 : NAND3_X1 port map( A1 => n354, A2 => n355, A3 => n226, ZN => n173);
   U310 : AOI22_X1 port map( A1 => A(15), A2 => n640, B1 => A(16), B2 => n630, 
                           ZN => n226);
   U311 : NAND3_X1 port map( A1 => n317, A2 => n318, A3 => n221, ZN => n168);
   U312 : AOI22_X1 port map( A1 => A(27), A2 => n639, B1 => A(28), B2 => n613, 
                           ZN => n221);
   U313 : OR2_X1 port map( A1 => n652, A2 => n621, ZN => n318);
   U314 : NAND2_X1 port map( A1 => SH(2), A2 => n228, ZN => n196);
   U315 : NAND2_X1 port map( A1 => n636, A2 => A(1), ZN => n350);
   U316 : OR2_X1 port map( A1 => n617, A2 => n682, ZN => n351);
   U317 : NAND3_X1 port map( A1 => n331, A2 => n332, A3 => n210, ZN => n166);
   U318 : AOI22_X1 port map( A1 => A(8), A2 => n639, B1 => A(9), B2 => n613, ZN
                           => n210);
   U319 : NAND2_X1 port map( A1 => n344, A2 => SH(0), ZN => n240);
   U320 : NOR2_X1 port map( A1 => n505, A2 => n506, ZN => n245);
   U321 : AND3_X1 port map( A1 => n362, A2 => n363, A3 => n364, ZN => n125);
   U322 : NAND2_X1 port map( A1 => n630, A2 => A(31), ZN => n362);
   U323 : NAND2_X1 port map( A1 => n639, A2 => A(30), ZN => n363);
   U324 : INV_X1 port map( A => A(31), ZN => n646);
   U325 : INV_X1 port map( A => A(23), ZN => n659);
   U326 : INV_X1 port map( A => A(6), ZN => n680);
   U327 : INV_X1 port map( A => A(28), ZN => n653);
   U328 : INV_X1 port map( A => A(26), ZN => n656);
   U329 : INV_X1 port map( A => A(19), ZN => n664);
   U330 : INV_X1 port map( A => A(17), ZN => n666);
   U331 : INV_X1 port map( A => A(16), ZN => n667);
   U332 : INV_X1 port map( A => A(9), ZN => n676);
   U333 : INV_X1 port map( A => A(22), ZN => n661);
   U334 : INV_X1 port map( A => A(13), ZN => n671);
   U335 : INV_X1 port map( A => A(18), ZN => n665);
   U336 : INV_X1 port map( A => A(20), ZN => n663);
   U337 : INV_X1 port map( A => A(25), ZN => n657);
   U338 : INV_X1 port map( A => A(5), ZN => n681);
   U339 : INV_X1 port map( A => A(27), ZN => n654);
   U340 : INV_X1 port map( A => A(30), ZN => n650);
   U341 : INV_X1 port map( A => A(8), ZN => n677);
   U342 : INV_X1 port map( A => A(7), ZN => n678);
   U343 : INV_X1 port map( A => A(21), ZN => n662);
   U344 : INV_X1 port map( A => A(24), ZN => n658);
   U345 : INV_X1 port map( A => A(14), ZN => n670);
   U346 : INV_X1 port map( A => A(12), ZN => n672);
   U347 : INV_X1 port map( A => A(11), ZN => n673);
   U348 : INV_X1 port map( A => A(0), ZN => n689);
   U349 : INV_X1 port map( A => A(15), ZN => n669);
   U350 : INV_X1 port map( A => A(29), ZN => n652);
   U351 : INV_X1 port map( A => A(3), ZN => n684);
   U352 : AND3_X1 port map( A1 => n248, A2 => SH(27), A3 => n309, ZN => n243);
   U353 : OAI22_X1 port map( A1 => n688, A2 => n104, B1 => n107, B2 => n181, ZN
                           => B(1));
   U354 : NAND2_X1 port map( A1 => n154, A2 => n625, ZN => n489);
   U355 : NAND2_X1 port map( A1 => n154, A2 => n642, ZN => n482);
   U356 : INV_X1 port map( A => A(2), ZN => n685);
   U357 : AOI22_X1 port map( A1 => A(2), A2 => n638, B1 => A(3), B2 => n613, ZN
                           => n197);
   U358 : AOI22_X1 port map( A1 => A(4), A2 => n639, B1 => A(5), B2 => n632, ZN
                           => n212);
   U359 : AOI22_X1 port map( A1 => A(3), A2 => n640, B1 => A(4), B2 => n632, ZN
                           => n220);
   U360 : INV_X1 port map( A => A(4), ZN => n682);
   U361 : AOI22_X1 port map( A1 => A(10), A2 => n640, B1 => A(11), B2 => n631, 
                           ZN => n199);
   U362 : AOI22_X1 port map( A1 => A(9), A2 => n640, B1 => A(10), B2 => n632, 
                           ZN => n232);
   U363 : INV_X1 port map( A => A(10), ZN => n675);
   U364 : OAI221_X1 port map( B1 => n594, B2 => n689, C1 => n620, C2 => n684, A
                           => n231, ZN => n153);
   U365 : AOI22_X1 port map( A1 => A(1), A2 => n639, B1 => A(2), B2 => n631, ZN
                           => n231);
   U366 : NAND2_X1 port map( A1 => n604, A2 => n584, ZN => n616);
   U367 : INV_X1 port map( A => n637, ZN => n635);
   U368 : OAI221_X1 port map( B1 => n133, B2 => n692, C1 => n134, C2 => n693, A
                           => n135, ZN => B(27));
   U369 : OAI22_X1 port map( A1 => n189, A2 => n690, B1 => n190, B2 => n693, ZN
                           => B(16));
   U370 : OAI22_X1 port map( A1 => n645, A2 => n112, B1 => n113, B2 => n114, ZN
                           => B(31));
   U371 : INV_X1 port map( A => n624, ZN => n617);
   U372 : INV_X1 port map( A => n599, ZN => n618);
   U374 : INV_X1 port map( A => n624, ZN => n619);
   U375 : INV_X1 port map( A => n597, ZN => n620);
   U376 : INV_X1 port map( A => n597, ZN => n621);
   U377 : INV_X1 port map( A => n599, ZN => n622);
   U378 : INV_X1 port map( A => n598, ZN => n623);
   U379 : NOR3_X1 port map( A1 => n329, A2 => n330, A3 => n660, ZN => n92);
   U380 : INV_X1 port map( A => n572, ZN => n683);
   U381 : AOI22_X1 port map( A1 => n587, A2 => n628, B1 => n572, B2 => n642, ZN
                           => n91);
   U382 : NAND2_X1 port map( A1 => n636, A2 => A(29), ZN => n364);
   U383 : NAND4_X1 port map( A1 => n244, A2 => n243, A3 => n245, A4 => n610, ZN
                           => n283);
   U384 : NAND4_X1 port map( A1 => n242, A2 => n244, A3 => n245, A4 => n243, ZN
                           => n241);
   U385 : AND3_X1 port map( A1 => SH(18), A2 => SH(17), A3 => SH(19), ZN => 
                           n247);
   U386 : NAND2_X1 port map( A1 => n241, A2 => SH(31), ZN => n344);
   U387 : NAND2_X1 port map( A1 => SH(31), A2 => n283, ZN => n228);
   U388 : INV_X1 port map( A => SH(31), ZN => n694);
   U389 : AND2_X1 port map( A1 => n136, A2 => n696, ZN => n376);
   U390 : NOR2_X1 port map( A1 => n196, A2 => n696, ZN => n387);
   U391 : NOR2_X1 port map( A1 => n697, A2 => n137, ZN => n261);
   U392 : INV_X1 port map( A => n137, ZN => n696);
   U393 : AOI222_X1 port map( A1 => n600, A2 => n643, B1 => n686, B2 => n626, 
                           C1 => n586, C2 => n628, ZN => n133);
   U394 : AOI22_X1 port map( A1 => n600, A2 => n633, B1 => n629, B2 => n592, ZN
                           => n184);
   U395 : AOI22_X1 port map( A1 => n598, A2 => A(1), B1 => n632, B2 => A(0), ZN
                           => n121);
   U396 : NOR2_X1 port map( A1 => n604, A2 => n383, ZN => n272);
   U397 : INV_X1 port map( A => n383, ZN => n698);
   U398 : AOI22_X1 port map( A1 => n633, A2 => n603, B1 => n629, B2 => n145, ZN
                           => n188);
   U399 : AOI222_X1 port map( A1 => n603, A2 => n643, B1 => n627, B2 => n143, 
                           C1 => n144, C2 => n628, ZN => n88);
   U400 : OAI222_X1 port map( A1 => n388, A2 => n690, B1 => n645, B2 => n191, 
                           C1 => n352, C2 => n693, ZN => B(15));
   U401 : OR2_X1 port map( A1 => n616, A2 => n662, ZN => n290);
   U402 : OR2_X1 port map( A1 => n635, A2 => n682, ZN => n294);
   U403 : OR2_X1 port map( A1 => n596, A2 => n676, ZN => n305);
   U404 : OR2_X1 port map( A1 => n616, A2 => n677, ZN => n314);
   U405 : OR2_X1 port map( A1 => n596, A2 => n658, ZN => n367);
   U406 : OR2_X1 port map( A1 => n594, A2 => n657, ZN => n371);
   U407 : OR2_X1 port map( A1 => n616, A2 => n663, ZN => n302);
   U408 : OR2_X1 port map( A1 => n616, A2 => n681, ZN => n286);
   U409 : OR2_X1 port map( A1 => n596, A2 => n684, ZN => n279);
   U410 : OR2_X1 port map( A1 => n594, A2 => n656, ZN => n317);
   U411 : OR2_X1 port map( A1 => n594, A2 => n673, ZN => n379);
   U412 : OR2_X1 port map( A1 => n596, A2 => n664, ZN => n365);
   U413 : OR2_X1 port map( A1 => n616, A2 => n672, ZN => n335);
   U414 : OR2_X1 port map( A1 => n596, A2 => n654, ZN => n342);
   U415 : OR2_X1 port map( A1 => n594, A2 => n669, ZN => n358);
   U416 : AOI22_X1 port map( A1 => n634, A2 => n173, B1 => n629, B2 => n168, ZN
                           => n195);
   U417 : OAI22_X1 port map( A1 => n117, A2 => n112, B1 => n113, B2 => n118, ZN
                           => B(30));
   U418 : OR2_X1 port map( A1 => n618, A2 => n666, ZN => n355);
   U419 : OR2_X1 port map( A1 => n616, A2 => n670, ZN => n354);
   U420 : OAI222_X1 port map( A1 => n127, A2 => n690, B1 => n125, B2 => n191, 
                           C1 => n322, C2 => n693, ZN => B(13));
   U421 : AOI222_X1 port map( A1 => n148, A2 => n629, B1 => n144, B2 => n642, 
                           C1 => n137, C2 => n101, ZN => n322);
   U422 : OR3_X1 port map( A1 => SH(14), A2 => SH(15), A3 => SH(13), ZN => n258
                           );
   U423 : OR2_X1 port map( A1 => n596, A2 => n678, ZN => n331);
   U424 : OR2_X1 port map( A1 => n621, A2 => n675, ZN => n332);
   U425 : NOR4_X1 port map( A1 => n257, A2 => SH(16), A3 => SH(18), A4 => n593,
                           ZN => n252);
   U426 : OR3_X1 port map( A1 => SH(20), A2 => SH(21), A3 => SH(19), ZN => n257
                           );
   U427 : OR3_X1 port map( A1 => SH(26), A2 => SH(27), A3 => SH(25), ZN => n256
                           );
   U428 : OAI221_X1 port map( B1 => n134, B2 => n690, C1 => n133, C2 => n693, A
                           => n208, ZN => B(11));
   U429 : INV_X1 port map( A => n213, ZN => n655);
   U430 : AND3_X1 port map( A1 => SH(24), A2 => SH(23), A3 => SH(25), ZN => 
                           n248);
   U431 : NOR4_X1 port map( A1 => n258, A2 => SH(10), A3 => SH(12), A4 => 
                           SH(11), ZN => n251);
   U432 : NAND4_X1 port map( A1 => SH(10), A2 => SH(12), A3 => SH(11), A4 => 
                           SH(13), ZN => n505);
   U433 : OR4_X1 port map( A1 => SH(6), A2 => SH(7), A3 => SH(8), A4 => SH(9), 
                           ZN => n255);
   U434 : AND3_X1 port map( A1 => SH(30), A2 => SH(29), A3 => SH(6), ZN => n249
                           );
   U435 : NOR4_X1 port map( A1 => n255, A2 => n611, A3 => SH(30), A4 => SH(29),
                           ZN => n254);
   U436 : AND2_X1 port map( A1 => SH(28), A2 => SH(26), ZN => n309);
   U437 : AOI221_X1 port map( B1 => n167, B2 => n626, C1 => n583, C2 => n641, A
                           => n649, ZN => n388);
   U438 : AND2_X1 port map( A1 => n167, A2 => n627, ZN => n356);
   U439 : AND2_X1 port map( A1 => n167, A2 => n634, ZN => n374);
   U440 : AOI22_X1 port map( A1 => n634, A2 => n586, B1 => n629, B2 => n167, ZN
                           => n165);
   U441 : NOR4_X1 port map( A1 => n256, A2 => SH(22), A3 => SH(24), A4 => 
                           SH(23), ZN => n253);
   U442 : INV_X1 port map( A => n615, ZN => n629);
   U443 : INV_X1 port map( A => n595, ZN => n636);
   U444 : INV_X1 port map( A => n595, ZN => n637);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity SHIFTER_M32_N5_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (31 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_M32_N5_DW01_ash_0;

architecture SYN_mx2 of SHIFTER_M32_N5_DW01_ash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal temp_int_SH_4_port, SHMAG_5_port, MR_int_1_31_port, MR_int_1_30_port,
      MR_int_1_29_port, MR_int_1_28_port, MR_int_1_27_port, MR_int_1_26_port, 
      MR_int_1_25_port, MR_int_1_24_port, MR_int_1_22_port, MR_int_1_21_port, 
      MR_int_1_16_port, MR_int_1_15_port, MR_int_1_14_port, MR_int_1_13_port, 
      MR_int_1_12_port, MR_int_1_11_port, MR_int_1_10_port, MR_int_1_9_port, 
      MR_int_1_8_port, MR_int_1_7_port, MR_int_1_6_port, MR_int_1_5_port, 
      MR_int_1_4_port, MR_int_1_3_port, MR_int_1_2_port, MR_int_1_1_port, 
      MR_int_2_31_port, MR_int_2_30_port, MR_int_2_29_port, MR_int_2_27_port, 
      MR_int_2_26_port, MR_int_2_25_port, MR_int_2_24_port, MR_int_2_23_port, 
      MR_int_2_22_port, MR_int_2_21_port, MR_int_2_20_port, MR_int_2_19_port, 
      MR_int_2_16_port, MR_int_2_15_port, MR_int_2_11_port, MR_int_2_10_port, 
      MR_int_2_9_port, MR_int_2_8_port, MR_int_2_7_port, MR_int_2_6_port, 
      MR_int_2_5_port, MR_int_2_4_port, MR_int_2_3_port, MR_int_2_2_port, 
      MR_int_2_1_port, MR_int_3_31_port, MR_int_3_30_port, MR_int_3_29_port, 
      MR_int_3_27_port, MR_int_3_26_port, MR_int_3_25_port, MR_int_3_24_port, 
      MR_int_3_23_port, MR_int_3_21_port, MR_int_3_20_port, MR_int_3_19_port, 
      MR_int_3_18_port, MR_int_3_17_port, MR_int_3_16_port, MR_int_3_15_port, 
      MR_int_3_12_port, MR_int_3_11_port, MR_int_3_10_port, MR_int_3_9_port, 
      MR_int_3_8_port, MR_int_3_7_port, MR_int_3_6_port, MR_int_3_4_port, 
      MR_int_3_3_port, MR_int_3_2_port, MR_int_3_1_port, MR_int_4_31_port, 
      MR_int_4_29_port, MR_int_4_28_port, MR_int_4_25_port, MR_int_4_24_port, 
      MR_int_4_22_port, MR_int_4_20_port, MR_int_4_19_port, MR_int_4_18_port, 
      MR_int_4_13_port, MR_int_4_12_port, MR_int_4_11_port, MR_int_4_10_port, 
      MR_int_4_8_port, MR_int_4_6_port, MR_int_4_4_port, MR_int_4_3_port, 
      MR_int_4_2_port, MR_int_5_3_port, MR_int_7_30_port, MR_int_7_29_port, 
      MR_int_7_24_port, MR_int_7_22_port, MR_int_7_20_port, MR_int_7_16_port, 
      ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, ML_int_1_28_port, 
      ML_int_1_26_port, ML_int_1_25_port, ML_int_1_24_port, ML_int_1_23_port, 
      ML_int_1_22_port, ML_int_1_21_port, ML_int_1_19_port, ML_int_1_18_port, 
      ML_int_1_17_port, ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, 
      ML_int_1_13_port, ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, 
      ML_int_1_9_port, ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, 
      ML_int_1_5_port, ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, 
      ML_int_1_1_port, ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, 
      ML_int_2_29_port, ML_int_2_28_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_21_port, ML_int_2_20_port, 
      ML_int_2_19_port, ML_int_2_17_port, ML_int_2_16_port, ML_int_2_15_port, 
      ML_int_2_14_port, ML_int_2_13_port, ML_int_2_12_port, ML_int_2_11_port, 
      ML_int_2_10_port, ML_int_2_9_port, ML_int_2_8_port, ML_int_2_7_port, 
      ML_int_2_6_port, ML_int_2_5_port, ML_int_2_4_port, ML_int_2_3_port, 
      ML_int_2_2_port, ML_int_2_1_port, ML_int_2_0_port, ML_int_3_31_port, 
      ML_int_3_30_port, ML_int_3_29_port, ML_int_3_28_port, ML_int_3_27_port, 
      ML_int_3_26_port, ML_int_3_25_port, ML_int_3_24_port, ML_int_3_23_port, 
      ML_int_3_21_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, ML_int_3_8_port, 
      ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, ML_int_3_4_port, 
      ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, ML_int_3_0_port, 
      ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, ML_int_4_28_port, 
      ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, ML_int_4_24_port, 
      ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, ML_int_4_20_port, 
      ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, ML_int_4_15_port, 
      ML_int_4_14_port, ML_int_4_13_port, ML_int_4_12_port, ML_int_4_11_port, 
      ML_int_4_10_port, ML_int_4_9_port, ML_int_4_8_port, ML_int_5_31_port, 
      ML_int_5_30_port, ML_int_5_26_port, ML_int_5_25_port, ML_int_5_24_port, 
      ML_int_5_23_port, ML_int_5_22_port, ML_int_5_21_port, ML_int_5_20_port, 
      ML_int_5_18_port, ML_int_5_17_port, ML_int_7_29_port, ML_int_7_28_port, 
      ML_int_7_16_port, ML_int_7_14_port, ML_int_7_10_port, ML_int_7_9_port, 
      ML_int_7_7_port, ML_int_7_6_port, ML_int_7_5_port, ML_int_7_3_port, 
      ML_int_7_2_port, ML_int_7_1_port, ML_int_7_0_port, n15, n80, n81, n82, 
      n84, n85, n86, n87, n88, n90, n92, n98, n104, net60450, net60477, 
      net60578, net60604, net60660, net60751, net60750, net60763, net60869, 
      net60893, net61039, net61046, net61053, net61132, net61266, net61331, 
      net61353, net61364, net61363, net61624, net61724, net61755, net61774, 
      net61783, net61782, net61842, net61851, ML_int_1_20_port, 
      ML_int_3_22_port, ML_int_2_22_port, ML_int_2_18_port, net65464, net65465,
      temp_int_SH_0_port, net61465, n99, n97, n91, n101, n100, MR_int_2_14_port
      , MR_int_4_30_port, MR_int_1_20_port, MR_int_1_18_port, net60718, 
      ML_int_7_13_port, net61436, net60589, net60588, MR_int_4_14_port, 
      MR_int_3_22_port, MR_int_3_14_port, MR_int_2_18_port, n121, n122, n124, 
      n125, n131, n132, n135, n136, n138, n139, n141, n142, n144, n145, n147, 
      n148, n150, n151, n153, n154, n155, n156, n157, n158, n160, n161, n162, 
      n163, n164, n168, n170, n171, n173, n174, n175, n178, n180, n181, n182, 
      n183, n184, n186, n189, n192, n193, n195, n196, n197, n199, n200, n201, 
      n204, n205, n207, n208, n210, n211, n212, n213, n214, n215, n219, n220, 
      n221, n223, n224, n225, n226, n227, n228, n229, n230, n232, n233, n234, 
      n235, n236, n237, n241, n243, n244, n245, n246, n250, n251, n252, n253, 
      n255, n256, n257, n261, n264, n267, n270, n271, n272, n273, n274, n279, 
      n282, n283, n284, n285, n286, n295, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
      n315, n318, n319, n320, n321, n324, n325, n326, n327, n328, n329, n331, 
      n332, n333, n334, n335, n336, n337, n338, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n369, n370, 
      n375, n376, n377, n378, n379, n380, n381, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n502, n503, n505, n506, n507, n508, n509, n510, n511, n512, 
      n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, 
      n525, n526, n527, n528, n529, n530, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n549, n550, n551, 
      n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
      n564, n565, n566, n567, n568, n569, n570, n571, n572, n574, n575, n576, 
      n577, n578, n579, n580, n581, n583, n584, n585, n586, n587, n588, n589, 
      n590, n591, n592, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n622, n623, n624, 
      n627, n628, net131991, net134827, net134825, net134821, net134819, 
      net134815, net134813, net134811, net134809, net134837, net134833, 
      net134831, net134867, net134865, net134861, net134859, net134855, 
      net134853, net134851, net134849, net134847, net134845, net134843, 
      net134839, net134881, net134879, net134875, net134913, net134911, 
      net134905, net134903, net134901, net134899, net134897, net134895, 
      net134893, net134891, net134889, net134887, net134885, net134883, 
      net134929, net134927, net134925, net134923, net134967, net134963, 
      net134959, net134957, net134953, net134951, net134949, net134947, 
      net134945, net134943, net134941, net134939, net134937, net134935, 
      net134933, net134971, net134969, net134977, net134975, net135715, 
      net135717, net135729, net135734, net135859, net135858, net135867, 
      net135866, net135876, net135875, net141178, net141255, net141408, 
      net141430, net141429, net141428, net141444, net141464, net141501, 
      net141507, net141516, net141528, net141534, net141544, net141543, 
      net141562, net141563, net141573, n290, n289, n288, n287, n109, n108, n107
      , n106, n96, n89, MR_int_1_19_port, net60313, n292, n291, n110, 
      temp_int_SH_3_port, temp_int_SH_1_port, net60576, net141212, net135865, 
      n95, MR_int_1_17_port, temp_int_SH_2_port, net134965, net134909, n548, 
      n547, n260, MR_int_2_17_port, MR_int_2_13_port, net135874, net131988, n83
      , n340, ML_int_7_4_port, net134961, net134873, net134863, 
      MR_int_3_13_port, net134871, net134869, net134841, n128, n127, 
      MR_int_4_5_port, MR_int_3_5_port, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
      n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
      n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, 
      n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
      n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, 
      n758 : std_logic;

begin
   
   M1_3_3 : MUX2_X1 port map( A => MR_int_3_3_port, B => MR_int_3_11_port, S =>
                           net134837, Z => MR_int_4_3_port);
   M1_3_2 : MUX2_X1 port map( A => MR_int_3_2_port, B => MR_int_3_10_port, S =>
                           net134831, Z => MR_int_4_2_port);
   M1_2_6_0 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_10_port, S 
                           => net134929, Z => MR_int_3_6_port);
   M1_2_4_0 : MUX2_X1 port map( A => MR_int_2_4_port, B => MR_int_2_8_port, S 
                           => net134927, Z => MR_int_3_4_port);
   M1_2_3 : MUX2_X1 port map( A => MR_int_2_3_port, B => MR_int_2_7_port, S => 
                           net134929, Z => MR_int_3_3_port);
   M1_1_11_0 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_13_port, 
                           S => net135859, Z => MR_int_2_11_port);
   M1_1_10_0 : MUX2_X1 port map( A => MR_int_1_10_port, B => MR_int_1_12_port, 
                           S => net135858, Z => MR_int_2_10_port);
   M1_1_4_0 : MUX2_X1 port map( A => MR_int_1_4_port, B => MR_int_1_6_port, S 
                           => net141464, Z => MR_int_2_4_port);
   M1_1_3_0 : MUX2_X1 port map( A => MR_int_1_3_port, B => MR_int_1_5_port, S 
                           => net135859, Z => MR_int_2_3_port);
   M1_1_1 : MUX2_X1 port map( A => MR_int_1_1_port, B => ML_int_1_4_port, S => 
                           net141464, Z => MR_int_2_1_port);
   M1_0_29_0 : MUX2_X1 port map( A => A(29), B => A(30), S => net141563, Z => 
                           MR_int_1_29_port);
   M1_0_28_0 : MUX2_X1 port map( A => A(28), B => A(29), S => net141408, Z => 
                           MR_int_1_28_port);
   M1_0_24_0 : MUX2_X1 port map( A => A(24), B => A(25), S => net131991, Z => 
                           MR_int_1_24_port);
   M1_0_22_0 : MUX2_X1 port map( A => A(22), B => A(23), S => net141516, Z => 
                           MR_int_1_22_port);
   M1_0_9_0 : MUX2_X1 port map( A => A(9), B => A(10), S => n742, Z => 
                           MR_int_1_9_port);
   M1_0_8_0 : MUX2_X1 port map( A => A(8), B => A(9), S => n742, Z => 
                           MR_int_1_8_port);
   M1_0_6_0 : MUX2_X1 port map( A => A(6), B => A(7), S => net135729, Z => 
                           MR_int_1_6_port);
   M1_0_5_0 : MUX2_X1 port map( A => A(5), B => A(6), S => net141255, Z => 
                           MR_int_1_5_port);
   M1_0_4_0 : MUX2_X1 port map( A => A(4), B => A(5), S => n695, Z => 
                           MR_int_1_4_port);
   M1_0_2_0 : MUX2_X1 port map( A => A(2), B => A(3), S => net141516, Z => 
                           MR_int_1_2_port);
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => net134811, Z => ML_int_5_25_port);
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => n755, S => net134811
                           , Z => ML_int_5_18_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => net134855, Z => ML_int_4_21_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => net134905, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => net134903, Z => ML_int_2_30_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => n297, S => net134903
                           , Z => ML_int_2_28_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           net134901, Z => ML_int_2_3_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n693, Z => 
                           ML_int_1_31_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n693, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => net141430, Z => 
                           ML_int_1_28_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => net141428, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => net141429, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => net61851, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => net61851, Z => 
                           ML_int_1_23_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n705, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n693, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => net141429, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => net135865, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n705, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => net135865, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => net61851, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => net141428, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n710, Z => 
                           ML_int_1_8_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => net135866, Z => 
                           ML_int_1_5_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => net135865, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => net61851, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => net141430, Z => 
                           ML_int_1_1_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => net141428, Z => 
                           ML_int_1_7_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => net141430, Z => 
                           ML_int_1_4_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => net141430, Z => 
                           ML_int_1_6_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => net134905, Z => ML_int_2_24_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n694, Z => 
                           ML_int_1_22_port);
   M1_0_13_0 : MUX2_X1 port map( A => A(13), B => A(14), S => n742, Z => 
                           MR_int_1_13_port);
   M1_0_1_0 : MUX2_X1 port map( A => A(1), B => A(2), S => net135729, Z => 
                           MR_int_1_1_port);
   M1_3_22_0 : MUX2_X1 port map( A => n727, B => MR_int_3_30_port, S => 
                           net134837, Z => MR_int_4_22_port);
   M1_3_11_0 : MUX2_X1 port map( A => MR_int_3_11_port, B => MR_int_3_19_port, 
                           S => net134837, Z => MR_int_4_11_port);
   M1_3_14_0 : MUX2_X1 port map( A => n669, B => n727, S => net134833, Z => 
                           MR_int_4_14_port);
   M1_2_27_0 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, 
                           S => net134923, Z => MR_int_3_27_port);
   U3 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_30_port, S => 
                           net134923, Z => ML_int_3_30_port);
   U9 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_2_port, S => 
                           net134953, Z => MR_int_3_2_port);
   U47 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_31_port, S => 
                           net134833, Z => ML_int_4_31_port);
   U78 : MUX2_X1 port map( A => ML_int_7_16_port, B => MR_int_7_16_port, S => 
                           net135876, Z => B(16));
   U93 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S => 
                           net134855, Z => ML_int_4_22_port);
   U127 : MUX2_X1 port map( A => A(22), B => A(23), S => net141534, Z => n186);
   U197 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, S => 
                           net134923, Z => n236);
   U204 : MUX2_X1 port map( A => MR_int_3_10_port, B => MR_int_3_18_port, S => 
                           net134837, Z => MR_int_4_10_port);
   U226 : MUX2_X1 port map( A => MR_int_2_11_port, B => MR_int_2_7_port, S => 
                           net134953, Z => MR_int_3_7_port);
   U228 : MUX2_X1 port map( A => MR_int_1_9_port, B => MR_int_1_7_port, S => 
                           net134905, Z => MR_int_2_7_port);
   U235 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S => 
                           net134903, Z => ML_int_2_13_port);
   U236 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_22_port, S => 
                           net134927, Z => ML_int_3_22_port);
   U241 : MUX2_X1 port map( A => ML_int_1_11_port, B => n728, S => net134881, Z
                           => n264);
   U248 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_17_port, S => 
                           net134833, Z => ML_int_4_17_port);
   U254 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_26_port, S => 
                           n692, Z => ML_int_2_26_port);
   U269 : NAND3_X1 port map( A1 => ML_int_5_25_port, A2 => n85, A3 => net134977
                           , ZN => n336);
   U271 : NAND3_X1 port map( A1 => ML_int_5_24_port, A2 => n85, A3 => net134977
                           , ZN => n527);
   U288 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_18_port, S => 
                           net134903, Z => MR_int_2_18_port);
   U294 : MUX2_X1 port map( A => MR_int_3_22_port, B => MR_int_3_30_port, S => 
                           net134831, Z => net61774);
   U370 : MUX2_X1 port map( A => MR_int_3_4_port, B => MR_int_3_12_port, S => 
                           net134837, Z => MR_int_4_4_port);
   U374 : MUX2_X1 port map( A => A(26), B => A(25), S => n705, Z => n297);
   U389 : MUX2_X1 port map( A => A(11), B => A(10), S => n693, Z => 
                           MR_int_1_10_port);
   U448 : MUX2_X1 port map( A => A(8), B => A(7), S => net141430, Z => 
                           MR_int_1_7_port);
   U493 : MUX2_X1 port map( A => A(28), B => A(27), S => n710, Z => 
                           MR_int_1_27_port);
   U557 : MUX2_X1 port map( A => A(4), B => A(3), S => n693, Z => 
                           MR_int_1_3_port);
   U558 : MUX2_X1 port map( A => A(30), B => A(31), S => net141212, Z => 
                           MR_int_1_30_port);
   U565 : MUX2_X1 port map( A => A(13), B => A(12), S => net141429, Z => 
                           MR_int_1_12_port);
   U601 : MUX2_X1 port map( A => MR_int_1_12_port, B => MR_int_1_14_port, S => 
                           net135858, Z => n410);
   U621 : MUX2_X1 port map( A => A(27), B => A(26), S => net141429, Z => n424);
   U734 : MUX2_X1 port map( A => A(16), B => A(15), S => n694, Z => 
                           MR_int_1_15_port);
   U768 : MUX2_X1 port map( A => A(15), B => A(14), S => n729, Z => 
                           MR_int_1_14_port);
   U777 : MUX2_X1 port map( A => MR_int_3_16_port, B => MR_int_3_8_port, S => 
                           net134855, Z => MR_int_4_8_port);
   U913 : MUX2_X1 port map( A => A(23), B => A(24), S => n742, Z => n601);
   U299 : MUX2_X1 port map( A => n424, B => ML_int_1_25_port, S => net134901, Z
                           => n250);
   U732 : MUX2_X1 port map( A => ML_int_7_29_port, B => MR_int_7_29_port, S => 
                           net135876, Z => B(29));
   U273 : AND2_X2 port map( A1 => SHMAG_5_port, A2 => net134977, ZN => n85);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           net134953, Z => ML_int_3_4_port);
   U365 : NAND3_X1 port map( A1 => SH(16), A2 => SH(15), A3 => SH(14), ZN => 
                           net60751);
   U364 : NAND3_X1 port map( A1 => SH(18), A2 => SH(17), A3 => SH(19), ZN => 
                           net61363);
   U281 : NAND3_X1 port map( A1 => SH(22), A2 => SH(21), A3 => SH(20), ZN => 
                           net61364);
   M1_0_20_0 : MUX2_X1 port map( A => A(20), B => A(21), S => net141408, Z => 
                           MR_int_1_20_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => net61851, Z => 
                           ML_int_1_20_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n710, Z => 
                           ML_int_1_21_port);
   U367 : NAND3_X1 port map( A1 => SH(8), A2 => SH(7), A3 => SH(9), ZN => 
                           net65464);
   U368 : NAND3_X1 port map( A1 => SH(30), A2 => SH(29), A3 => SH(6), ZN => 
                           net65465);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => net61851, Z => 
                           ML_int_1_19_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => net141429, Z => 
                           ML_int_1_17_port);
   M1_0_16_0 : MUX2_X1 port map( A => A(16), B => A(17), S => net141563, Z => 
                           MR_int_1_16_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => net141544, Z => 
                           ML_int_1_18_port);
   M1_0_25_0 : MUX2_X1 port map( A => A(25), B => A(26), S => net141212, Z => 
                           MR_int_1_25_port);
   M1_0_17_0 : MUX2_X1 port map( A => A(17), B => A(18), S => net141178, Z => 
                           MR_int_1_17_port);
   M1_2_5_0 : MUX2_X1 port map( A => MR_int_2_5_port, B => MR_int_2_9_port, S 
                           => net134925, Z => MR_int_3_5_port);
   U4 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n107, A4 => n108, ZN 
                           => n656);
   U5 : BUF_X1 port map( A => temp_int_SH_0_port, Z => net135865);
   U6 : AND3_X1 port map( A1 => n657, A2 => n658, A3 => n659, ZN => n109);
   U7 : NOR2_X1 port map( A1 => SH(27), A2 => SH(26), ZN => n657);
   U8 : AND2_X1 port map( A1 => n721, A2 => n719, ZN => n658);
   U10 : AND2_X1 port map( A1 => n720, A2 => n718, ZN => n659);
   U11 : BUF_X1 port map( A => net134961, Z => net134939);
   U12 : NAND2_X1 port map( A1 => MR_int_3_26_port, A2 => net134833, ZN => n660
                           );
   U13 : INV_X1 port map( A => net141501, ZN => net141429);
   U14 : INV_X2 port map( A => net134967, ZN => net134925);
   U15 : NAND2_X1 port map( A1 => MR_int_3_17_port, A2 => n664, ZN => n661);
   U16 : NAND2_X1 port map( A1 => n661, A2 => n662, ZN => MR_int_7_16_port);
   U17 : OR2_X1 port map( A1 => n663, A2 => n243, ZN => n662);
   U18 : INV_X1 port map( A => n205, ZN => n663);
   U19 : AND2_X1 port map( A1 => net134839, A2 => n205, ZN => n664);
   U20 : CLKBUF_X1 port map( A => n579, Z => n665);
   U21 : BUF_X2 port map( A => net134911, Z => net134897);
   U22 : NAND2_X1 port map( A1 => n723, A2 => n666, ZN => B(11));
   U23 : AND2_X1 port map( A1 => n724, A2 => n532, ZN => n666);
   U24 : INV_X2 port map( A => net141501, ZN => net141430);
   U25 : NAND2_X1 port map( A1 => MR_int_4_14_port, A2 => n170, ZN => n667);
   U26 : NAND2_X1 port map( A1 => n667, A2 => n668, ZN => B(13));
   U27 : AND2_X1 port map( A1 => net60718, A2 => n168, ZN => n668);
   U28 : NAND2_X1 port map( A1 => net60588, A2 => net60589, ZN => n669);
   U29 : MUX2_X1 port map( A => A(30), B => A(29), S => net135867, Z => 
                           ML_int_1_30_port);
   U30 : CLKBUF_X1 port map( A => n689, Z => n670);
   U31 : BUF_X1 port map( A => temp_int_SH_2_port, Z => net134967);
   U32 : INV_X1 port map( A => net134965, ZN => net134929);
   U33 : BUF_X1 port map( A => net134911, Z => net134883);
   U34 : INV_X1 port map( A => temp_int_SH_2_port, ZN => net134927);
   U35 : INV_X1 port map( A => net134827, ZN => net134811);
   U36 : BUF_X1 port map( A => net134911, Z => net134903);
   U37 : NAND2_X1 port map( A1 => net134927, A2 => net134865, ZN => n671);
   U38 : NAND2_X1 port map( A1 => n85, A2 => net134977, ZN => n672);
   U39 : NAND2_X1 port map( A1 => MR_int_3_1_port, A2 => net134855, ZN => n673)
                           ;
   U40 : BUF_X1 port map( A => SH(31), Z => net135875);
   U41 : BUF_X1 port map( A => net131988, Z => net134975);
   U42 : MUX2_X1 port map( A => MR_int_3_12_port, B => MR_int_3_20_port, S => 
                           net134837, Z => MR_int_4_12_port);
   U43 : CLKBUF_X1 port map( A => SH(31), Z => net135874);
   U44 : MUX2_X1 port map( A => MR_int_1_13_port, B => MR_int_1_15_port, S => 
                           net134881, Z => MR_int_2_13_port);
   U45 : BUF_X1 port map( A => temp_int_SH_1_port, Z => net134909);
   U46 : MUX2_X1 port map( A => A(19), B => A(18), S => net141544, Z => 
                           MR_int_1_18_port);
   U48 : BUF_X1 port map( A => SH(31), Z => net135876);
   U49 : AND2_X1 port map( A1 => n303, A2 => n304, ZN => n674);
   U50 : NOR2_X1 port map( A1 => n675, A2 => n676, ZN => n679);
   U51 : AND2_X1 port map( A1 => n606, A2 => n607, ZN => n675);
   U52 : NAND2_X1 port map( A1 => net134971, A2 => n716, ZN => n676);
   U53 : OAI21_X1 port map( B1 => n678, B2 => n679, A => net135875, ZN => n677)
                           ;
   U54 : AND2_X1 port map( A1 => MR_int_4_5_port, A2 => n205, ZN => n678);
   U55 : OAI21_X1 port map( B1 => net134925, B2 => n680, A => n503, ZN => 
                           ML_int_3_19_port);
   U56 : INV_X1 port map( A => ML_int_2_15_port, ZN => n680);
   U57 : OAI221_X1 port map( B1 => n681, B2 => n476, C1 => n224, C2 => n737, A 
                           => n502, ZN => B(0));
   U58 : INV_X1 port map( A => n295, ZN => n681);
   U59 : AOI22_X1 port map( A1 => n731, A2 => ML_int_1_21_port, B1 => n682, B2 
                           => net134923, ZN => n510);
   U60 : INV_X1 port map( A => n459, ZN => n682);
   U61 : NAND3_X1 port map( A1 => n422, A2 => n225, A3 => n423, ZN => n163);
   U62 : NAND2_X1 port map( A1 => n344, A2 => n343, ZN => ML_int_2_15_port);
   U63 : OAI21_X1 port map( B1 => n683, B2 => n670, A => net134833, ZN => n468)
                           ;
   U64 : INV_X1 port map( A => n565, ZN => n683);
   U65 : OAI21_X1 port map( B1 => n674, B2 => n672, A => n572, ZN => B(19));
   U66 : OAI21_X1 port map( B1 => net134827, B2 => n673, A => n744, ZN => n295)
                           ;
   U67 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S => 
                           temp_int_SH_2_port, Z => ML_int_3_26_port);
   U68 : AOI21_X1 port map( B1 => n193, B2 => n192, A => net134825, ZN => n684)
                           ;
   U69 : INV_X1 port map( A => n684, ZN => n533);
   U70 : AOI21_X1 port map( B1 => n702, B2 => n701, A => n685, ZN => n686);
   U71 : INV_X1 port map( A => n493, ZN => n685);
   U72 : INV_X1 port map( A => n686, ZN => n402);
   U73 : NAND2_X1 port map( A1 => n299, A2 => n298, ZN => ML_int_5_26_port);
   U74 : NAND3_X1 port map( A1 => n232, A2 => n233, A3 => n594, ZN => B(9));
   U75 : NAND2_X1 port map( A1 => net134879, A2 => MR_int_1_14_port, ZN => n343
                           );
   U76 : INV_X2 port map( A => net134911, ZN => net134879);
   U77 : OAI22_X1 port map( A1 => n687, A2 => n671, B1 => net61039, B2 => 
                           net134837, ZN => n688);
   U79 : INV_X1 port map( A => n348, ZN => n687);
   U80 : INV_X1 port map( A => n688, ZN => n489);
   U81 : NAND3_X1 port map( A1 => n363, A2 => n409, A3 => n364, ZN => 
                           ML_int_4_9_port);
   U82 : AOI21_X1 port map( B1 => n547, B2 => n548, A => net134923, ZN => n689)
                           ;
   U83 : INV_X1 port map( A => n689, ZN => n564);
   U84 : AOI21_X1 port map( B1 => n468, B2 => n467, A => net134825, ZN => n690)
                           ;
   U85 : INV_X1 port map( A => n690, ZN => n411);
   U86 : AOI21_X1 port map( B1 => n589, B2 => n588, A => n476, ZN => n691);
   U87 : INV_X1 port map( A => n691, ZN => n610);
   U88 : INV_X1 port map( A => net134905, ZN => n692);
   U89 : BUF_X2 port map( A => net134909, Z => net134905);
   U90 : BUF_X1 port map( A => net135734, Z => n693);
   U91 : BUF_X1 port map( A => n729, Z => n694);
   U92 : BUF_X1 port map( A => temp_int_SH_0_port, Z => net141544);
   U94 : BUF_X1 port map( A => net134913, Z => net134901);
   U95 : BUF_X1 port map( A => net134967, Z => net134959);
   U96 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_18_port, S => 
                           net134897, Z => net61353);
   U97 : INV_X1 port map( A => net141544, ZN => n695);
   U98 : AND2_X1 port map( A1 => n583, A2 => n213, ZN => n696);
   U99 : NAND2_X1 port map( A1 => ML_int_4_22_port, A2 => net134815, ZN => n697
                           );
   U100 : NAND2_X1 port map( A1 => n752, A2 => net134811, ZN => n698);
   U101 : NAND2_X1 port map( A1 => n697, A2 => n698, ZN => ML_int_5_22_port);
   U102 : CLKBUF_X1 port map( A => net134913, Z => net134887);
   U103 : CLKBUF_X1 port map( A => net134911, Z => net134885);
   U104 : NAND2_X1 port map( A1 => ML_int_1_5_port, A2 => net135859, ZN => n699
                           );
   U105 : NAND2_X1 port map( A1 => ML_int_1_3_port, A2 => net134903, ZN => n700
                           );
   U106 : NAND2_X1 port map( A1 => n699, A2 => n700, ZN => ML_int_2_5_port);
   U107 : AND2_X2 port map( A1 => n96, A2 => n89, ZN => net141501);
   U108 : NAND2_X1 port map( A1 => ML_int_4_11_port, A2 => net134813, ZN => 
                           n701);
   U109 : NAND2_X1 port map( A1 => ML_int_4_27_port, A2 => net134815, ZN => 
                           n702);
   U110 : BUF_X1 port map( A => temp_int_SH_0_port, Z => net141543);
   U111 : NAND2_X1 port map( A1 => MR_int_4_24_port, A2 => net134811, ZN => 
                           n703);
   U112 : OR2_X1 port map( A1 => n703, A2 => n704, ZN => n515);
   U113 : OR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => n704);
   U114 : BUF_X1 port map( A => net135734, Z => n705);
   U115 : NAND2_X1 port map( A1 => MR_int_1_25_port, A2 => net134879, ZN => 
                           n706);
   U116 : NAND2_X1 port map( A1 => n601, A2 => net134903, ZN => n707);
   U117 : NAND2_X1 port map( A1 => n706, A2 => n707, ZN => MR_int_2_23_port);
   U118 : AND2_X1 port map( A1 => n708, A2 => n709, ZN => n446);
   U119 : NAND2_X1 port map( A1 => MR_int_4_13_port, A2 => n204, ZN => n708);
   U120 : OR2_X1 port map( A1 => n359, A2 => n456, ZN => n709);
   U121 : BUF_X1 port map( A => net135734, Z => n710);
   U122 : NAND2_X1 port map( A1 => ML_int_1_30_port, A2 => n711, ZN => n712);
   U123 : NAND2_X1 port map( A1 => MR_int_1_27_port, A2 => net134901, ZN => 
                           n713);
   U124 : NAND2_X1 port map( A1 => n712, A2 => n713, ZN => MR_int_2_27_port);
   U125 : INV_X1 port map( A => net134901, ZN => n711);
   U126 : NAND2_X1 port map( A1 => ML_int_4_30_port, A2 => net134815, ZN => 
                           n714);
   U128 : NAND2_X1 port map( A1 => ML_int_4_14_port, A2 => net134811, ZN => 
                           n715);
   U129 : NAND2_X1 port map( A1 => n714, A2 => n715, ZN => ML_int_5_30_port);
   U130 : INV_X1 port map( A => SHMAG_5_port, ZN => n716);
   U131 : AND2_X1 port map( A1 => net134813, A2 => n716, ZN => n205);
   U132 : NAND2_X1 port map( A1 => n716, A2 => n274, ZN => n271);
   U133 : BUF_X2 port map( A => n173, Z => net134971);
   U134 : NAND2_X1 port map( A1 => n127, A2 => n128, ZN => MR_int_4_5_port);
   U135 : NAND2_X1 port map( A1 => MR_int_3_5_port, A2 => net134841, ZN => n128
                           );
   U136 : BUF_X1 port map( A => net134869, Z => net134841);
   U137 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => net134841, ZN => n491
                           );
   U138 : NAND2_X1 port map( A1 => MR_int_3_21_port, A2 => net134841, ZN => 
                           n606);
   U139 : NAND2_X1 port map( A1 => ML_int_3_18_port, A2 => net134841, ZN => 
                           n145);
   U140 : BUF_X1 port map( A => net134871, Z => net134869);
   U141 : BUF_X1 port map( A => net134869, Z => net134839);
   U142 : BUF_X1 port map( A => net134869, Z => net134843);
   U143 : AND2_X1 port map( A1 => net134971, A2 => net134869, ZN => n220);
   U144 : CLKBUF_X1 port map( A => temp_int_SH_3_port, Z => net134871);
   U145 : CLKBUF_X1 port map( A => net134871, Z => net134867);
   U146 : INV_X1 port map( A => net134871, ZN => net134837);
   U147 : NAND2_X1 port map( A1 => MR_int_3_13_port, A2 => net134833, ZN => 
                           n127);
   U148 : INV_X2 port map( A => net134859, ZN => net134833);
   U149 : BUF_X2 port map( A => net134863, Z => net134859);
   U150 : BUF_X1 port map( A => net134873, Z => net134863);
   U151 : CLKBUF_X1 port map( A => net134863, Z => net134861);
   U152 : BUF_X1 port map( A => temp_int_SH_3_port, Z => net134873);
   U153 : BUF_X1 port map( A => net134873, Z => net134865);
   U154 : MUX2_X1 port map( A => MR_int_2_17_port, B => MR_int_2_13_port, S => 
                           net134939, Z => MR_int_3_13_port);
   U155 : BUF_X1 port map( A => net134965, Z => net134961);
   U156 : BUF_X1 port map( A => net134961, Z => net134941);
   U157 : BUF_X1 port map( A => net134961, Z => net134943);
   U158 : BUF_X1 port map( A => temp_int_SH_2_port, Z => net134965);
   U159 : NAND2_X1 port map( A1 => n677, A2 => n340, ZN => B(4));
   U160 : NAND2_X1 port map( A1 => ML_int_7_4_port, A2 => net134977, ZN => n340
                           );
   U161 : BUF_X4 port map( A => net131988, Z => net134977);
   U162 : INV_X1 port map( A => net135874, ZN => net131988);
   U163 : NAND2_X1 port map( A1 => n106, A2 => net131988, ZN => net61465);
   U164 : NAND2_X1 port map( A1 => n656, A2 => net131988, ZN => n89);
   U165 : NOR2_X1 port map( A1 => n325, A2 => n83, ZN => ML_int_7_4_port);
   U166 : NAND2_X1 port map( A1 => net141573, A2 => net134833, ZN => n83);
   U167 : BUF_X1 port map( A => net134965, Z => net134963);
   U168 : NAND2_X1 port map( A1 => n547, A2 => n548, ZN => MR_int_2_17_port);
   U169 : MUX2_X1 port map( A => MR_int_2_13_port, B => MR_int_2_17_port, S => 
                           net134929, Z => net141562);
   U170 : NAND2_X1 port map( A1 => MR_int_1_19_port, A2 => net134875, ZN => 
                           n548);
   U171 : INV_X1 port map( A => net134905, ZN => net134875);
   U172 : INV_X1 port map( A => net134909, ZN => net135717);
   U173 : NAND2_X1 port map( A1 => MR_int_1_17_port, A2 => net134897, ZN => 
                           n547);
   U174 : BUF_X2 port map( A => temp_int_SH_1_port, Z => net134911);
   U175 : NAND2_X1 port map( A1 => MR_int_2_13_port, A2 => net134927, ZN => 
                           n557);
   U176 : NAND2_X1 port map( A1 => net61465, A2 => n260, ZN => 
                           temp_int_SH_2_port);
   U177 : INV_X1 port map( A => temp_int_SH_2_port, ZN => net134923);
   U178 : NAND2_X1 port map( A1 => SH(2), A2 => net141507, ZN => n260);
   U179 : NAND2_X1 port map( A1 => MR_int_1_19_port, A2 => net134891, ZN => 
                           n595);
   U180 : CLKBUF_X1 port map( A => temp_int_SH_1_port, Z => net134913);
   U181 : NAND2_X1 port map( A1 => MR_int_1_17_port, A2 => net134879, ZN => 
                           n581);
   U182 : INV_X1 port map( A => net135867, ZN => net141212);
   U183 : INV_X1 port map( A => net135867, ZN => net131991);
   U184 : NAND2_X1 port map( A1 => n89, A2 => n95, ZN => temp_int_SH_1_port);
   U185 : NAND2_X1 port map( A1 => SH(1), A2 => net60576, ZN => n95);
   U186 : NAND2_X1 port map( A1 => net60578, A2 => net135875, ZN => net60576);
   U187 : NAND2_X1 port map( A1 => n89, A2 => n96, ZN => temp_int_SH_0_port);
   U188 : CLKBUF_X1 port map( A => net61465, Z => net135715);
   U189 : NAND2_X1 port map( A1 => net60578, A2 => net135875, ZN => net141507);
   U190 : NAND2_X1 port map( A1 => net61465, A2 => n717, ZN => 
                           temp_int_SH_3_port);
   U191 : NAND2_X1 port map( A1 => SH(3), A2 => net141507, ZN => n717);
   U192 : AND3_X1 port map( A1 => net60313, A2 => n292, A3 => n291, ZN => n110)
                           ;
   U193 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n107, A4 => n108, ZN
                           => n106);
   U194 : NOR2_X1 port map( A1 => SH(6), A2 => SH(9), ZN => n291);
   U195 : NOR2_X1 port map( A1 => SH(8), A2 => SH(7), ZN => n292);
   U196 : NOR3_X1 port map( A1 => SH(28), A2 => SH(29), A3 => SH(30), ZN => 
                           net60313);
   U198 : AND3_X1 port map( A1 => SH(28), A2 => SH(26), A3 => SH(27), ZN => 
                           net60450);
   U199 : MUX2_X1 port map( A => A(20), B => A(19), S => net141430, Z => 
                           MR_int_1_19_port);
   U200 : NAND2_X1 port map( A1 => n91, A2 => SH(0), ZN => n96);
   U201 : NAND2_X1 port map( A1 => n91, A2 => SH(0), ZN => net141444);
   U202 : AND2_X1 port map( A1 => n287, A2 => n289, ZN => n108);
   U203 : NOR3_X1 port map( A1 => SH(20), A2 => SH(21), A3 => SH(19), ZN => 
                           n289);
   U205 : NOR3_X1 port map( A1 => SH(17), A2 => SH(18), A3 => SH(16), ZN => 
                           n287);
   U206 : AND2_X1 port map( A1 => n290, A2 => n288, ZN => n107);
   U207 : NOR3_X1 port map( A1 => SH(11), A2 => SH(12), A3 => SH(10), ZN => 
                           n288);
   U208 : NOR3_X1 port map( A1 => SH(14), A2 => SH(15), A3 => SH(13), ZN => 
                           n290);
   U209 : INV_X1 port map( A => SH(22), ZN => n718);
   U210 : INV_X1 port map( A => SH(24), ZN => n720);
   U211 : INV_X1 port map( A => SH(23), ZN => n719);
   U212 : INV_X1 port map( A => SH(25), ZN => n721);
   U213 : NAND4_X1 port map( A1 => SH(11), A2 => SH(12), A3 => SH(13), A4 => 
                           SH(10), ZN => net60750);
   U214 : AND3_X1 port map( A1 => SH(24), A2 => SH(25), A3 => SH(23), ZN => 
                           n104);
   U215 : NAND2_X1 port map( A1 => ML_int_2_13_port, A2 => n722, ZN => n356);
   U216 : AND2_X1 port map( A1 => net134929, A2 => net134837, ZN => n722);
   U217 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           net134953, Z => net141573);
   U218 : NAND2_X1 port map( A1 => MR_int_4_12_port, A2 => n241, ZN => n723);
   U219 : OR2_X1 port map( A1 => n208, A2 => n592, ZN => n724);
   U220 : BUF_X1 port map( A => temp_int_SH_0_port, Z => net135866);
   U221 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, S => 
                           net134925, Z => n725);
   U222 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, S => 
                           net134923, Z => n726);
   U223 : NAND2_X1 port map( A1 => n279, A2 => net60477, ZN => n727);
   U224 : INV_X1 port map( A => net135866, ZN => net141563);
   U225 : MUX2_X1 port map( A => A(13), B => A(12), S => net141544, Z => n728);
   U227 : MUX2_X1 port map( A => A(27), B => A(26), S => net141429, Z => 
                           MR_int_1_26_port);
   U229 : INV_X1 port map( A => net141428, ZN => net141534);
   U230 : INV_X1 port map( A => net134905, ZN => net141528);
   U231 : INV_X1 port map( A => net141428, ZN => net141516);
   U232 : NAND2_X1 port map( A1 => net61465, A2 => net141444, ZN => n729);
   U233 : NAND2_X1 port map( A1 => net61465, A2 => net141444, ZN => net61851);
   U234 : INV_X1 port map( A => net134897, ZN => net141464);
   U237 : BUF_X2 port map( A => net135717, Z => net135858);
   U238 : INV_X1 port map( A => net141501, ZN => net141428);
   U239 : INV_X1 port map( A => net141543, ZN => net141408);
   U240 : NAND2_X1 port map( A1 => n484, A2 => n485, ZN => n730);
   U242 : AND2_X1 port map( A1 => net135858, A2 => net134927, ZN => n731);
   U243 : MUX2_X1 port map( A => A(12), B => A(11), S => net141430, Z => 
                           MR_int_1_11_port);
   U244 : MUX2_X1 port map( A => A(28), B => A(29), S => net141534, Z => n732);
   U245 : NAND2_X1 port map( A1 => ML_int_4_29_port, A2 => n733, ZN => n735);
   U246 : NOR2_X1 port map( A1 => n758, A2 => net134813, ZN => n733);
   U247 : MUX2_X2 port map( A => MR_int_2_30_port, B => MR_int_2_26_port, S => 
                           net134967, Z => MR_int_3_26_port);
   U249 : NAND2_X1 port map( A1 => ML_int_4_13_port, A2 => n736, ZN => n734);
   U250 : NAND2_X1 port map( A1 => n735, A2 => n734, ZN => ML_int_7_29_port);
   U251 : AND2_X1 port map( A1 => net134809, A2 => n85, ZN => n736);
   U252 : INV_X1 port map( A => net141543, ZN => net135729);
   U253 : INV_X1 port map( A => net135866, ZN => net141255);
   U255 : OR2_X1 port map( A1 => net134811, A2 => n476, ZN => n737);
   U256 : BUF_X2 port map( A => net134957, Z => net134953);
   U257 : BUF_X1 port map( A => net134957, Z => net134951);
   U258 : CLKBUF_X1 port map( A => net134911, Z => net134889);
   U259 : INV_X1 port map( A => net141543, ZN => net141178);
   U260 : INV_X1 port map( A => n88, ZN => n757);
   U261 : INV_X1 port map( A => n87, ZN => n756);
   U262 : NAND2_X1 port map( A1 => n753, A2 => net134809, ZN => n125);
   U263 : INV_X1 port map( A => n82, ZN => n753);
   U264 : OR2_X1 port map( A1 => net134811, A2 => n603, ZN => n183);
   U265 : INV_X1 port map( A => n84, ZN => n754);
   U266 : INV_X1 port map( A => net134825, ZN => net134809);
   U267 : AND2_X1 port map( A1 => n477, A2 => n256, ZN => n178);
   U268 : INV_X1 port map( A => net134905, ZN => net134881);
   U270 : NOR2_X1 port map( A1 => n325, A2 => n84, ZN => ML_int_7_3_port);
   U272 : NOR2_X1 port map( A1 => n325, A2 => n81, ZN => ML_int_7_6_port);
   U274 : BUF_X1 port map( A => net134865, Z => net134855);
   U275 : BUF_X1 port map( A => net134867, Z => net134847);
   U276 : NOR2_X1 port map( A1 => net134925, A2 => n751, ZN => MR_int_3_30_port
                           );
   U277 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => net134833, ZN => n84)
                           ;
   U278 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => net134833, ZN => n86)
                           ;
   U279 : CLKBUF_X1 port map( A => net134865, Z => net134853);
   U280 : BUF_X1 port map( A => net134963, Z => net134935);
   U282 : BUF_X1 port map( A => net134963, Z => net134933);
   U283 : BUF_X1 port map( A => net134867, Z => net134845);
   U284 : BUF_X1 port map( A => net134959, Z => net134945);
   U285 : BUF_X1 port map( A => net134867, Z => net134849);
   U286 : NAND2_X1 port map( A1 => ML_int_3_14_port, A2 => net134831, ZN => 
                           n550);
   U287 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => net134851, ZN => n551
                           );
   U289 : NAND2_X1 port map( A1 => n174, A2 => net134833, ZN => n423);
   U290 : NAND2_X1 port map( A1 => n445, A2 => n444, ZN => n174);
   U291 : BUF_X1 port map( A => net134865, Z => net134851);
   U292 : NAND2_X1 port map( A1 => n416, A2 => n415, ZN => ML_int_4_12_port);
   U293 : BUF_X1 port map( A => net134963, Z => net134937);
   U295 : BUF_X1 port map( A => net134959, Z => net134949);
   U296 : NAND2_X1 port map( A1 => n437, A2 => n438, ZN => ML_int_4_11_port);
   U297 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => net134847, ZN => n438
                           );
   U298 : NAND2_X1 port map( A1 => ML_int_3_11_port, A2 => net134837, ZN => 
                           n437);
   U300 : NAND2_X1 port map( A1 => n400, A2 => n399, ZN => ML_int_4_20_port);
   U301 : NAND2_X1 port map( A1 => n253, A2 => net134831, ZN => n399);
   U302 : NAND2_X1 port map( A1 => net61132, A2 => n475, ZN => ML_int_4_15_port
                           );
   U303 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => net134847, ZN => n475
                           );
   U304 : NAND2_X1 port map( A1 => ML_int_3_15_port, A2 => net134831, ZN => 
                           net61132);
   U305 : NAND2_X1 port map( A1 => ML_int_4_8_port, A2 => n622, ZN => n267);
   U306 : NAND2_X1 port map( A1 => n490, A2 => n491, ZN => ML_int_4_8_port);
   U307 : NAND2_X1 port map( A1 => ML_int_3_8_port, A2 => net134831, ZN => n490
                           );
   U308 : BUF_X1 port map( A => net134959, Z => net134947);
   U309 : NAND2_X1 port map( A1 => ML_int_3_16_port, A2 => net134853, ZN => 
                           n432);
   U310 : NAND2_X1 port map( A1 => ML_int_4_19_port, A2 => net134819, ZN => 
                           n303);
   U311 : NAND2_X1 port map( A1 => ML_int_3_11_port, A2 => net134845, ZN => 
                           n426);
   U312 : NAND2_X1 port map( A1 => n138, A2 => n139, ZN => ML_int_4_10_port);
   U313 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => net134847, ZN => n139
                           );
   U314 : NAND2_X1 port map( A1 => ML_int_5_17_port, A2 => n379, ZN => n450);
   U315 : NAND2_X1 port map( A1 => n360, A2 => n361, ZN => ML_int_5_17_port);
   U316 : NAND2_X1 port map( A1 => n756, A2 => net134809, ZN => n361);
   U317 : AND2_X1 port map( A1 => net134861, A2 => net134971, ZN => n184);
   U318 : NAND2_X1 port map( A1 => ML_int_5_20_port, A2 => n227, ZN => n443);
   U319 : NAND2_X1 port map( A1 => n366, A2 => n367, ZN => ML_int_5_20_port);
   U320 : NAND2_X1 port map( A1 => n309, A2 => net134809, ZN => n367);
   U321 : NAND2_X1 port map( A1 => ML_int_4_20_port, A2 => net134819, ZN => 
                           n366);
   U322 : NAND2_X1 port map( A1 => n513, A2 => n512, ZN => ML_int_4_23_port);
   U323 : NAND2_X1 port map( A1 => ML_int_3_23_port, A2 => net134831, ZN => 
                           n513);
   U324 : NAND2_X1 port map( A1 => ML_int_3_15_port, A2 => net134845, ZN => 
                           n512);
   U325 : NAND2_X1 port map( A1 => ML_int_3_22_port, A2 => net134847, ZN => 
                           net61053);
   U326 : AND2_X1 port map( A1 => ML_int_3_16_port, A2 => n158, ZN => n161);
   U327 : AND2_X1 port map( A1 => ML_int_3_8_port, A2 => n199, ZN => n160);
   U328 : AND2_X1 port map( A1 => net134861, A2 => n252, ZN => n199);
   U329 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n622, ZN => 
                           ML_int_7_9_port);
   U330 : NAND2_X1 port map( A1 => ML_int_3_8_port, A2 => n246, ZN => n244);
   U331 : OR2_X1 port map( A1 => n197, A2 => net134971, ZN => n388);
   U332 : OR2_X1 port map( A1 => n750, A2 => net134971, ZN => n324);
   U333 : INV_X1 port map( A => MR_int_4_28_port, ZN => n750);
   U334 : OR2_X1 port map( A1 => net134825, A2 => n491, ZN => n245);
   U335 : NAND2_X1 port map( A1 => ML_int_5_23_port, A2 => n379, ZN => n514);
   U336 : NAND2_X1 port map( A1 => n471, A2 => n472, ZN => ML_int_5_23_port);
   U337 : OR2_X1 port map( A1 => n80, A2 => net134827, ZN => n472);
   U338 : NAND2_X1 port map( A1 => ML_int_4_23_port, A2 => net134819, ZN => 
                           n471);
   U339 : OR2_X1 port map( A1 => n466, A2 => net134859, ZN => n364);
   U340 : NAND2_X1 port map( A1 => n470, A2 => n469, ZN => ML_int_5_24_port);
   U341 : NAND2_X1 port map( A1 => ML_int_4_24_port, A2 => net134969, ZN => 
                           n470);
   U342 : AND2_X1 port map( A1 => n244, A2 => n245, ZN => n469);
   U343 : NAND2_X1 port map( A1 => n431, A2 => n432, ZN => ML_int_4_24_port);
   U344 : INV_X1 port map( A => n86, ZN => n755);
   U345 : NAND2_X1 port map( A1 => n369, A2 => n370, ZN => ML_int_4_18_port);
   U346 : NAND2_X1 port map( A1 => n430, A2 => n429, ZN => ML_int_4_27_port);
   U347 : NAND2_X1 port map( A1 => n328, A2 => n329, ZN => ML_int_7_16_port);
   U348 : OR2_X1 port map( A1 => n758, A2 => n362, ZN => n329);
   U349 : NOR2_X1 port map( A1 => n160, A2 => n161, ZN => n328);
   U350 : NAND2_X1 port map( A1 => n757, A2 => net134811, ZN => n362);
   U351 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n622, ZN => 
                           ML_int_7_10_port);
   U352 : NAND2_X1 port map( A1 => ML_int_5_22_port, A2 => n493, ZN => n495);
   U353 : INV_X1 port map( A => n81, ZN => n752);
   U354 : INV_X1 port map( A => n225, ZN => n746);
   U355 : NAND2_X1 port map( A1 => n85, A2 => net134969, ZN => n325);
   U356 : AND2_X1 port map( A1 => n85, A2 => net134971, ZN => n622);
   U357 : NAND2_X1 port map( A1 => ML_int_7_9_port, A2 => net134975, ZN => n594
                           );
   U358 : NAND2_X1 port map( A1 => ML_int_4_11_port, A2 => n211, ZN => n532);
   U359 : NAND2_X1 port map( A1 => n455, A2 => n454, ZN => B(15));
   U360 : NAND2_X1 port map( A1 => n384, A2 => n622, ZN => n455);
   U361 : NAND2_X1 port map( A1 => n446, A2 => n447, ZN => B(12));
   U362 : NAND2_X1 port map( A1 => n235, A2 => n622, ZN => n447);
   U363 : BUF_X1 port map( A => n173, Z => net134969);
   U366 : AND2_X1 port map( A1 => ML_int_5_31_port, A2 => n378, ZN => B(31));
   U369 : AND2_X1 port map( A1 => n85, A2 => net134977, ZN => n378);
   U371 : AND2_X1 port map( A1 => net134813, A2 => n405, ZN => n383);
   U372 : NAND2_X1 port map( A1 => n402, A2 => n401, ZN => B(27));
   U373 : OR2_X1 port map( A1 => n324, A2 => n359, ZN => n401);
   U375 : NAND2_X1 port map( A1 => ML_int_7_13_port, A2 => net134975, ZN => 
                           net60718);
   U376 : NAND2_X1 port map( A1 => ML_int_2_6_port, A2 => net134927, ZN => n586
                           );
   U377 : NAND2_X1 port map( A1 => ML_int_2_2_port, A2 => net134941, ZN => n587
                           );
   U378 : AND2_X1 port map( A1 => net134977, A2 => n85, ZN => n493);
   U379 : NAND2_X1 port map( A1 => ML_int_7_5_port, A2 => net134975, ZN => n559
                           );
   U380 : NOR2_X1 port map( A1 => n82, A2 => n325, ZN => ML_int_7_5_port);
   U381 : NAND2_X1 port map( A1 => n433, A2 => n434, ZN => ML_int_3_8_port);
   U382 : NAND2_X1 port map( A1 => ML_int_2_8_port, A2 => net134927, ZN => n433
                           );
   U383 : NAND2_X1 port map( A1 => ML_int_2_4_port, A2 => net134943, ZN => n434
                           );
   U384 : NAND2_X1 port map( A1 => n171, A2 => net134833, ZN => n607);
   U385 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n622, ZN => 
                           ML_int_7_14_port);
   U386 : CLKBUF_X1 port map( A => net134913, Z => net134893);
   U387 : NAND2_X1 port map( A1 => MR_int_2_21_port, A2 => net134937, ZN => 
                           n478);
   U388 : NAND2_X1 port map( A1 => ML_int_2_6_port, A2 => net134939, ZN => n540
                           );
   U390 : NAND2_X1 port map( A1 => ML_int_2_12_port, A2 => net134927, ZN => 
                           n320);
   U391 : NAND2_X1 port map( A1 => ML_int_2_14_port, A2 => net134939, ZN => 
                           n521);
   U392 : NAND2_X1 port map( A1 => ML_int_2_18_port, A2 => net134927, ZN => 
                           net60893);
   U393 : NAND2_X1 port map( A1 => ML_int_2_5_port, A2 => net134925, ZN => n300
                           );
   U394 : AND2_X1 port map( A1 => n85, A2 => net134977, ZN => n227);
   U395 : AND2_X1 port map( A1 => n85, A2 => net134977, ZN => n379);
   U396 : NAND2_X1 port map( A1 => n507, A2 => n506, ZN => n253);
   U397 : NAND2_X1 port map( A1 => ML_int_2_20_port, A2 => net134927, ZN => 
                           n506);
   U398 : NAND2_X1 port map( A1 => n141, A2 => n142, ZN => ML_int_3_15_port);
   U399 : NAND2_X1 port map( A1 => ML_int_2_15_port, A2 => net134925, ZN => 
                           n141);
   U400 : NAND2_X1 port map( A1 => n538, A2 => n537, ZN => ML_int_3_11_port);
   U401 : NAND2_X1 port map( A1 => ML_int_2_7_port, A2 => net134941, ZN => n538
                           );
   U402 : CLKBUF_X1 port map( A => net134913, Z => net134891);
   U403 : CLKBUF_X1 port map( A => net134911, Z => net134899);
   U404 : AND2_X1 port map( A1 => net134827, A2 => n85, ZN => n252);
   U405 : OR2_X1 port map( A1 => n271, A2 => net134977, ZN => n335);
   U406 : NAND2_X1 port map( A1 => n345, A2 => n357, ZN => n355);
   U407 : NAND2_X1 port map( A1 => MR_int_2_23_port, A2 => net134923, ZN => 
                           n545);
   U408 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => net134925, ZN => 
                           ML_int_3_3_port);
   U409 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => net134925, ZN => 
                           ML_int_3_2_port);
   U410 : NAND2_X1 port map( A1 => ML_int_2_5_port, A2 => net134933, ZN => n466
                           );
   U411 : NAND2_X1 port map( A1 => n517, A2 => n516, ZN => ML_int_3_13_port);
   U412 : AND2_X1 port map( A1 => MR_int_3_29_port, A2 => net134843, ZN => 
                           MR_int_4_29_port);
   U413 : AND2_X1 port map( A1 => n623, A2 => n624, ZN => MR_int_4_28_port);
   U414 : INV_X1 port map( A => n85, ZN => n758);
   U415 : CLKBUF_X1 port map( A => net134911, Z => net134895);
   U416 : NAND2_X1 port map( A1 => n220, A2 => n221, ZN => n225);
   U417 : NOR2_X1 port map( A1 => n392, A2 => n162, ZN => n221);
   U418 : NAND2_X1 port map( A1 => net134953, A2 => net61436, ZN => n162);
   U419 : NAND2_X1 port map( A1 => ML_int_3_27_port, A2 => net134833, ZN => 
                           n430);
   U420 : NAND2_X1 port map( A1 => n480, A2 => n481, ZN => ML_int_3_27_port);
   U421 : NAND2_X1 port map( A1 => n250, A2 => net134923, ZN => n480);
   U422 : NAND2_X1 port map( A1 => ML_int_2_23_port, A2 => net134951, ZN => 
                           n481);
   U423 : NAND2_X1 port map( A1 => net61755, A2 => n349, ZN => MR_int_4_6_port)
                           ;
   U424 : NAND2_X1 port map( A1 => MR_int_3_6_port, A2 => net134849, ZN => n349
                           );
   U425 : NAND2_X1 port map( A1 => MR_int_3_14_port, A2 => net134831, ZN => 
                           net61755);
   U426 : NAND2_X1 port map( A1 => ML_int_3_24_port, A2 => net134837, ZN => 
                           n431);
   U427 : NAND2_X1 port map( A1 => n341, A2 => n342, ZN => ML_int_3_24_port);
   U428 : NAND2_X1 port map( A1 => ML_int_2_20_port, A2 => net134933, ZN => 
                           n342);
   U429 : NAND2_X1 port map( A1 => n518, A2 => n519, ZN => ML_int_3_16_port);
   U430 : NAND2_X1 port map( A1 => ML_int_2_12_port, A2 => net134945, ZN => 
                           n519);
   U431 : NAND2_X1 port map( A1 => n410, A2 => net134927, ZN => n407);
   U432 : NAND2_X1 port map( A1 => n484, A2 => n485, ZN => MR_int_3_24_port);
   U433 : NAND2_X1 port map( A1 => n473, A2 => n474, ZN => ML_int_3_7_port);
   U434 : NAND2_X1 port map( A1 => ML_int_2_3_port, A2 => net134943, ZN => n474
                           );
   U435 : NAND2_X1 port map( A1 => ML_int_2_7_port, A2 => net134925, ZN => n473
                           );
   U436 : NOR2_X1 port map( A1 => n325, A2 => n88, ZN => ML_int_7_0_port);
   U437 : NOR2_X1 port map( A1 => n325, A2 => n86, ZN => ML_int_7_2_port);
   U438 : NOR2_X1 port map( A1 => n325, A2 => n87, ZN => ML_int_7_1_port);
   U439 : NOR2_X1 port map( A1 => n80, A2 => n325, ZN => ML_int_7_7_port);
   U440 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => net134923, ZN => 
                           ML_int_3_0_port);
   U441 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => net134925, ZN => 
                           ML_int_3_1_port);
   U442 : NAND2_X1 port map( A1 => n375, A2 => n376, ZN => ML_int_7_28_port);
   U443 : NAND2_X1 port map( A1 => ML_int_4_28_port, A2 => n252, ZN => n376);
   U444 : NAND2_X1 port map( A1 => ML_int_4_12_port, A2 => n377, ZN => n375);
   U445 : NAND2_X1 port map( A1 => n552, A2 => n553, ZN => ML_int_3_14_port);
   U446 : NAND2_X1 port map( A1 => ML_int_2_14_port, A2 => net134923, ZN => 
                           n552);
   U447 : NAND2_X1 port map( A1 => n489, A2 => n488, ZN => ML_int_4_25_port);
   U449 : NAND2_X1 port map( A1 => ML_int_3_25_port, A2 => net134831, ZN => 
                           n488);
   U450 : NAND2_X1 port map( A1 => n466, A2 => n465, ZN => ML_int_3_9_port);
   U451 : NAND2_X1 port map( A1 => ML_int_3_29_port, A2 => net134831, ZN => 
                           n387);
   U452 : NAND2_X1 port map( A1 => MR_int_2_8_port, A2 => net134935, ZN => n406
                           );
   U453 : NAND2_X1 port map( A1 => ML_int_2_24_port, A2 => net134935, ZN => 
                           n418);
   U454 : AND2_X1 port map( A1 => net134811, A2 => n85, ZN => n377);
   U455 : AND2_X1 port map( A1 => net134811, A2 => n261, ZN => n234);
   U456 : NAND2_X1 port map( A1 => MR_int_3_18_port, A2 => net134839, ZN => 
                           n575);
   U457 : NAND2_X1 port map( A1 => n460, A2 => n461, ZN => B(6));
   U458 : NAND2_X1 port map( A1 => MR_int_4_22_port, A2 => n189, ZN => n428);
   U459 : NOR2_X1 port map( A1 => net134971, A2 => net61266, ZN => n189);
   U460 : OR2_X1 port map( A1 => n476, A2 => n180, ZN => n168);
   U461 : NAND2_X1 port map( A1 => MR_int_4_30_port, A2 => net134969, ZN => 
                           n180);
   U462 : NAND2_X1 port map( A1 => n754, A2 => net134809, ZN => n304);
   U463 : NAND2_X1 port map( A1 => n486, A2 => n487, ZN => ML_int_3_25_port);
   U464 : NAND2_X1 port map( A1 => ML_int_2_25_port, A2 => net134923, ZN => 
                           n486);
   U465 : NAND2_X1 port map( A1 => ML_int_5_26_port, A2 => n493, ZN => n525);
   U466 : NAND2_X1 port map( A1 => ML_int_4_26_port, A2 => net134821, ZN => 
                           n298);
   U467 : NAND2_X1 port map( A1 => n163, A2 => n164, ZN => n568);
   U468 : OR2_X1 port map( A1 => n746, A2 => n226, ZN => n164);
   U469 : AND2_X1 port map( A1 => net134811, A2 => n306, ZN => n226);
   U470 : NAND2_X1 port map( A1 => n450, A2 => n451, ZN => B(17));
   U471 : OR2_X1 port map( A1 => n210, A2 => n541, ZN => n451);
   U472 : NAND2_X1 port map( A1 => n525, A2 => n524, ZN => B(26));
   U473 : OR2_X1 port map( A1 => n388, A2 => net60660, ZN => n524);
   U474 : NAND2_X1 port map( A1 => n156, A2 => n157, ZN => n572);
   U475 : NOR2_X1 port map( A1 => net134969, A2 => net60660, ZN => n157);
   U476 : NAND2_X1 port map( A1 => n427, A2 => n428, ZN => B(21));
   U477 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => net134853, ZN => n409
                           );
   U478 : NAND2_X1 port map( A1 => n345, A2 => n365, ZN => n363);
   U479 : NAND2_X1 port map( A1 => n181, A2 => net61436, ZN => n558);
   U480 : NAND2_X1 port map( A1 => ML_int_5_21_port, A2 => net61624, ZN => n427
                           );
   U481 : AND2_X1 port map( A1 => n85, A2 => net134977, ZN => net61624);
   U482 : NAND2_X1 port map( A1 => n124, A2 => n125, ZN => ML_int_5_21_port);
   U483 : NAND2_X1 port map( A1 => ML_int_4_21_port, A2 => net134821, ZN => 
                           n124);
   U484 : AND2_X1 port map( A1 => n622, A2 => net134977, ZN => n211);
   U485 : AND2_X1 port map( A1 => net134813, A2 => n237, ZN => n204);
   U486 : AND2_X1 port map( A1 => net134813, A2 => n405, ZN => n241);
   U487 : OR2_X1 port map( A1 => n358, A2 => n359, ZN => n435);
   U488 : NAND2_X1 port map( A1 => n223, A2 => net134809, ZN => n358);
   U489 : NAND2_X1 port map( A1 => n738, A2 => n739, ZN => n454);
   U490 : NAND2_X1 port map( A1 => n627, A2 => n628, ZN => n738);
   U491 : NOR2_X1 port map( A1 => net134971, A2 => net61266, ZN => n739);
   U492 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => net134977, ZN => n384
                           );
   U494 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => net134977, ZN => n235
                           );
   U495 : NAND2_X1 port map( A1 => n272, A2 => n273, ZN => n499);
   U496 : NAND2_X1 port map( A1 => MR_int_4_25_port, A2 => net134969, ZN => 
                           n412);
   U497 : NAND2_X1 port map( A1 => n308, A2 => n307, ZN => MR_int_3_12_port);
   U498 : NAND2_X1 port map( A1 => n410, A2 => net134951, ZN => n307);
   U499 : NAND2_X1 port map( A1 => net61331, A2 => n439, ZN => MR_int_3_10_port
                           );
   U500 : NAND2_X1 port map( A1 => MR_int_2_10_port, A2 => net134953, ZN => 
                           n439);
   U501 : NAND2_X1 port map( A1 => n131, A2 => n132, ZN => ML_int_5_31_port);
   U502 : NAND2_X1 port map( A1 => ML_int_4_31_port, A2 => net134815, ZN => 
                           n131);
   U503 : NAND2_X1 port map( A1 => ML_int_4_15_port, A2 => net134809, ZN => 
                           n132);
   U504 : AND2_X1 port map( A1 => net134971, A2 => n549, ZN => n201);
   U505 : NAND2_X1 port map( A1 => MR_int_4_28_port, A2 => net134969, ZN => 
                           n592);
   U506 : NAND2_X1 port map( A1 => ML_int_2_25_port, A2 => net134949, ZN => 
                           n390);
   U507 : NAND2_X1 port map( A1 => ML_int_5_30_port, A2 => n421, ZN => n529);
   U508 : AND2_X1 port map( A1 => n85, A2 => net134977, ZN => n421);
   U509 : AND2_X1 port map( A1 => net134811, A2 => n273, ZN => n214);
   U510 : AND2_X1 port map( A1 => net134811, A2 => net61436, ZN => n170);
   U511 : NAND2_X1 port map( A1 => MR_int_3_16_port, A2 => net134853, ZN => 
                           n627);
   U512 : OR2_X1 port map( A1 => net60660, A2 => net134971, ZN => n210);
   U513 : OR2_X1 port map( A1 => n359, A2 => n449, ZN => n256);
   U514 : AND2_X1 port map( A1 => net134859, A2 => net134971, ZN => n175);
   U515 : OR2_X1 port map( A1 => n207, A2 => n208, ZN => n319);
   U516 : OR2_X1 port map( A1 => n748, A2 => net134971, ZN => n207);
   U517 : INV_X1 port map( A => MR_int_4_29_port, ZN => n748);
   U518 : NAND2_X1 port map( A1 => MR_int_4_8_port, A2 => n257, ZN => n255);
   U519 : AND2_X1 port map( A1 => net134811, A2 => n237, ZN => n257);
   U520 : NAND2_X1 port map( A1 => n406, A2 => n407, ZN => MR_int_3_8_port);
   U521 : NAND2_X1 port map( A1 => n229, A2 => n230, ZN => n233);
   U522 : NAND2_X1 port map( A1 => MR_int_4_10_port, A2 => n234, ZN => n232);
   U523 : AND2_X1 port map( A1 => n237, A2 => net134971, ZN => n230);
   U524 : NAND2_X1 port map( A1 => MR_int_4_29_port, A2 => net134969, ZN => 
                           n456);
   U525 : NOR2_X1 port map( A1 => SHMAG_5_port, A2 => net134975, ZN => net61436
                           );
   U526 : NOR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => n237);
   U527 : AND2_X1 port map( A1 => n602, A2 => n603, ZN => n580);
   U528 : NOR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => n273);
   U529 : NOR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => n405);
   U530 : NOR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => n549);
   U531 : NOR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => n261);
   U532 : NAND2_X1 port map( A1 => n696, A2 => n212, ZN => B(3));
   U533 : NOR2_X1 port map( A1 => SHMAG_5_port, A2 => net134975, ZN => n306);
   U534 : NAND2_X1 port map( A1 => ML_int_1_18_port, A2 => net134891, ZN => 
                           net61783);
   U535 : NAND2_X1 port map( A1 => ML_int_1_10_port, A2 => net134885, ZN => 
                           n483);
   U536 : NAND2_X1 port map( A1 => ML_int_1_5_port, A2 => net134885, ZN => n441
                           );
   U537 : NAND2_X1 port map( A1 => ML_int_1_6_port, A2 => net134885, ZN => n492
                           );
   U538 : NOR2_X1 port map( A1 => net134971, A2 => SHMAG_5_port, ZN => n391);
   U539 : AND2_X1 port map( A1 => MR_int_4_25_port, A2 => n391, ZN => 
                           MR_int_7_24_port);
   U540 : NAND2_X1 port map( A1 => ML_int_1_19_port, A2 => net134893, ZN => 
                           n459);
   U541 : NAND2_X1 port map( A1 => MR_int_1_7_port, A2 => net134893, ZN => n398
                           );
   U542 : NAND2_X1 port map( A1 => MR_int_1_14_port, A2 => net134887, ZN => 
                           n282);
   U543 : NAND2_X1 port map( A1 => ML_int_1_16_port, A2 => net134889, ZN => 
                           net60604);
   U544 : NAND2_X1 port map( A1 => n200, A2 => n505, ZN => ML_int_2_9_port);
   U545 : OR2_X1 port map( A1 => net134977, A2 => SHMAG_5_port, ZN => n359);
   U546 : NAND2_X1 port map( A1 => n728, A2 => net134887, ZN => n344);
   U547 : NAND2_X1 port map( A1 => n508, A2 => n509, ZN => ML_int_2_14_port);
   U548 : NAND2_X1 port map( A1 => ML_int_1_12_port, A2 => net134887, ZN => 
                           n509);
   U549 : NAND2_X1 port map( A1 => n452, A2 => n453, ZN => ML_int_2_25_port);
   U550 : NAND2_X1 port map( A1 => ML_int_1_23_port, A2 => net134887, ZN => 
                           n453);
   U551 : NAND2_X1 port map( A1 => n393, A2 => n394, ZN => ML_int_2_6_port);
   U552 : NAND2_X1 port map( A1 => MR_int_1_3_port, A2 => net134889, ZN => n394
                           );
   U553 : NAND2_X1 port map( A1 => ML_int_2_17_port, A2 => net134945, ZN => 
                           n511);
   U554 : NAND2_X1 port map( A1 => n457, A2 => n302, ZN => ML_int_2_17_port);
   U555 : OR2_X1 port map( A1 => net134977, A2 => SHMAG_5_port, ZN => net60660)
                           ;
   U556 : NAND2_X1 port map( A1 => ML_int_1_7_port, A2 => net134883, ZN => n505
                           );
   U559 : NAND2_X1 port map( A1 => n530, A2 => net60869, ZN => ML_int_2_4_port)
                           ;
   U560 : NAND2_X1 port map( A1 => ML_int_1_2_port, A2 => net134897, ZN => n530
                           );
   U561 : NAND2_X1 port map( A1 => n608, A2 => n609, ZN => MR_int_2_21_port);
   U562 : NAND2_X1 port map( A1 => MR_int_1_21_port, A2 => net134891, ZN => 
                           n608);
   U563 : NAND2_X1 port map( A1 => n195, A2 => n196, ZN => ML_int_2_2_port);
   U564 : NAND2_X1 port map( A1 => ML_int_1_0_port, A2 => net134893, ZN => n196
                           );
   U566 : NAND2_X1 port map( A1 => n121, A2 => n122, ZN => ML_int_2_23_port);
   U567 : NAND2_X1 port map( A1 => ML_int_1_21_port, A2 => net134885, ZN => 
                           n122);
   U568 : NOR2_X1 port map( A1 => SHMAG_5_port, A2 => n15, ZN => 
                           MR_int_7_29_port);
   U569 : OR2_X1 port map( A1 => net134971, A2 => n743, ZN => n15);
   U570 : NAND2_X1 port map( A1 => n497, A2 => n498, ZN => MR_int_2_8_port);
   U571 : NAND2_X1 port map( A1 => MR_int_1_8_port, A2 => net134897, ZN => n497
                           );
   U572 : NAND2_X1 port map( A1 => n591, A2 => n590, ZN => MR_int_3_16_port);
   U573 : NAND2_X1 port map( A1 => net60588, A2 => net60589, ZN => 
                           MR_int_3_14_port);
   U574 : OR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => net61266)
                           ;
   U575 : NAND2_X1 port map( A1 => n326, A2 => n327, ZN => ML_int_2_18_port);
   U576 : NAND2_X1 port map( A1 => MR_int_1_15_port, A2 => net134895, ZN => 
                           n327);
   U577 : NAND2_X1 port map( A1 => ML_int_2_29_port, A2 => net134923, ZN => 
                           n389);
   U578 : NAND2_X1 port map( A1 => n413, A2 => n414, ZN => ML_int_2_29_port);
   U579 : NAND2_X1 port map( A1 => n424, A2 => net134883, ZN => n413);
   U580 : NAND2_X1 port map( A1 => n457, A2 => n302, ZN => n348);
   U581 : NAND2_X1 port map( A1 => n595, A2 => n596, ZN => MR_int_2_19_port);
   U582 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_9_port, S => 
                           net134903, Z => MR_int_2_9_port);
   U583 : OR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => n208);
   U584 : NAND2_X1 port map( A1 => ML_int_1_17_port, A2 => net134883, ZN => 
                           n353);
   U585 : NAND2_X1 port map( A1 => n568, A2 => n569, ZN => B(14));
   U586 : NAND2_X1 port map( A1 => n420, A2 => n419, ZN => ML_int_4_28_port);
   U587 : NAND2_X1 port map( A1 => ML_int_3_28_port, A2 => net134831, ZN => 
                           n419);
   U588 : NAND2_X1 port map( A1 => n253, A2 => net134849, ZN => n420);
   U589 : NAND2_X1 port map( A1 => n418, A2 => n417, ZN => ML_int_3_28_port);
   U590 : NAND2_X1 port map( A1 => n443, A2 => n442, ZN => B(20));
   U591 : NOR2_X1 port map( A1 => net134975, A2 => SHMAG_5_port, ZN => n313);
   U592 : AND2_X1 port map( A1 => n182, A2 => n183, ZN => n534);
   U593 : NAND2_X1 port map( A1 => n436, A2 => n435, ZN => B(18));
   U594 : NAND2_X1 port map( A1 => ML_int_5_18_port, A2 => n227, ZN => n436);
   U595 : AND2_X1 port map( A1 => MR_int_4_31_port, A2 => n391, ZN => 
                           MR_int_7_30_port);
   U596 : AND2_X1 port map( A1 => n598, A2 => n597, ZN => n305);
   U597 : INV_X1 port map( A => MR_int_1_31_port, ZN => n747);
   U598 : OR2_X1 port map( A1 => SHMAG_5_port, A2 => net134977, ZN => n476);
   U599 : NAND2_X1 port map( A1 => n311, A2 => n310, ZN => ML_int_2_22_port);
   U600 : NAND2_X1 port map( A1 => ML_int_1_20_port, A2 => net134897, ZN => 
                           n310);
   U602 : NAND2_X1 port map( A1 => n150, A2 => n151, ZN => ML_int_3_31_port);
   U603 : NAND2_X1 port map( A1 => n250, A2 => net134935, ZN => n150);
   U604 : NOR2_X1 port map( A1 => n740, A2 => n741, ZN => MR_int_7_20_port);
   U605 : AND2_X1 port map( A1 => n606, A2 => n607, ZN => n740);
   U606 : OR2_X1 port map( A1 => SHMAG_5_port, A2 => net134969, ZN => n741);
   U607 : INV_X1 port map( A => A(31), ZN => n749);
   U608 : MUX2_X1 port map( A => A(22), B => A(21), S => n705, Z => 
                           MR_int_1_21_port);
   U609 : NAND2_X1 port map( A1 => ML_int_1_15_port, A2 => net134899, ZN => 
                           n302);
   U610 : NAND2_X1 port map( A1 => MR_int_1_22_port, A2 => net134901, ZN => 
                           n561);
   U611 : NAND2_X1 port map( A1 => ML_int_2_28_port, A2 => net134923, ZN => 
                           n417);
   U612 : NAND2_X1 port map( A1 => MR_int_1_2_port, A2 => net134899, ZN => n154
                           );
   U613 : NAND2_X1 port map( A1 => n610, A2 => n611, ZN => B(1));
   U614 : NAND2_X1 port map( A1 => ML_int_3_30_port, A2 => net134837, ZN => 
                           n494);
   U615 : AND2_X1 port map( A1 => net134925, A2 => net134837, ZN => n365);
   U616 : AND2_X1 port map( A1 => net134837, A2 => n252, ZN => n158);
   U617 : AND2_X1 port map( A1 => net134837, A2 => net134811, ZN => n246);
   U618 : NAND2_X1 port map( A1 => n499, A2 => n500, ZN => B(8));
   U619 : BUF_X1 port map( A => temp_int_SH_0_port, Z => net135867);
   U620 : CLKBUF_X3 port map( A => net135717, Z => net135859);
   U622 : NAND2_X1 port map( A1 => SH(4), A2 => net141507, ZN => n90);
   U623 : NAND2_X1 port map( A1 => SH(5), A2 => net141507, ZN => n92);
   U624 : NOR2_X1 port map( A1 => net141464, A2 => n747, ZN => MR_int_2_31_port
                           );
   U625 : OR2_X1 port map( A1 => net135859, A2 => n747, ZN => n392);
   U626 : NAND2_X1 port map( A1 => MR_int_1_31_port, A2 => net135859, ZN => 
                           n598);
   U627 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => net135859, ZN => 
                           ML_int_2_0_port);
   U628 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => net135859, ZN => 
                           ML_int_2_1_port);
   U629 : NAND2_X1 port map( A1 => n228, A2 => net134833, ZN => n523);
   U630 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => net134831, ZN => n80)
                           ;
   U631 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => net134837, ZN => n87)
                           ;
   U632 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => net134837, ZN => n88)
                           ;
   U633 : NAND2_X1 port map( A1 => ML_int_1_9_port, A2 => net134879, ZN => n200
                           );
   U634 : NAND2_X1 port map( A1 => ML_int_1_17_port, A2 => net134879, ZN => 
                           n457);
   U635 : NAND2_X1 port map( A1 => ML_int_1_29_port, A2 => net134879, ZN => 
                           n414);
   U636 : NAND2_X1 port map( A1 => ML_int_1_25_port, A2 => net134879, ZN => 
                           n452);
   U637 : NAND2_X1 port map( A1 => net61465, A2 => net141444, ZN => net135734);
   U638 : INV_X1 port map( A => n729, ZN => n742);
   U639 : NAND2_X1 port map( A1 => n312, A2 => n313, ZN => n460);
   U640 : NAND2_X1 port map( A1 => MR_int_3_31_port, A2 => net134833, ZN => 
                           n603);
   U641 : AND2_X1 port map( A1 => net134861, A2 => MR_int_3_31_port, ZN => 
                           MR_int_4_31_port);
   U642 : NOR2_X1 port map( A1 => net134927, A2 => n392, ZN => MR_int_3_31_port
                           );
   U643 : NOR2_X1 port map( A1 => net134929, A2 => n215, ZN => n228);
   U644 : NOR2_X1 port map( A1 => net134929, A2 => n305, ZN => MR_int_3_29_port
                           );
   U645 : NOR2_X1 port map( A1 => net134929, A2 => n305, ZN => n171);
   U646 : NOR2_X1 port map( A1 => net134837, A2 => net134929, ZN => n624);
   U647 : NAND2_X1 port map( A1 => n348, A2 => net134929, ZN => n496);
   U648 : NAND2_X1 port map( A1 => ML_int_2_24_port, A2 => net134929, ZN => 
                           n341);
   U649 : NAND2_X1 port map( A1 => ML_int_2_31_port, A2 => net134929, ZN => 
                           n151);
   U650 : NAND2_X1 port map( A1 => ML_int_2_13_port, A2 => net134929, ZN => 
                           n516);
   U651 : AND2_X1 port map( A1 => net134963, A2 => net134837, ZN => n357);
   U652 : NAND2_X1 port map( A1 => n337, A2 => n338, ZN => MR_int_4_13_port);
   U653 : NAND2_X1 port map( A1 => net141562, A2 => net134853, ZN => n337);
   U654 : NAND2_X1 port map( A1 => n623, A2 => net134927, ZN => n484);
   U655 : NAND2_X1 port map( A1 => n251, A2 => net134845, ZN => n400);
   U656 : NAND2_X1 port map( A1 => n251, A2 => net134831, ZN => n415);
   U657 : NAND2_X1 port map( A1 => n492, A2 => n334, ZN => ML_int_2_8_port);
   U658 : BUF_X1 port map( A => net134967, Z => net134957);
   U659 : NAND2_X1 port map( A1 => n440, A2 => n441, ZN => ML_int_2_7_port);
   U660 : NAND2_X1 port map( A1 => ML_int_1_7_port, A2 => net141528, ZN => n440
                           );
   U661 : NAND2_X1 port map( A1 => MR_int_2_18_port, A2 => net134923, ZN => 
                           net60588);
   U662 : NAND2_X1 port map( A1 => n566, A2 => n567, ZN => MR_int_3_20_port);
   U663 : NAND2_X1 port map( A1 => MR_int_1_24_port, A2 => net134893, ZN => 
                           n599);
   U664 : NAND2_X1 port map( A1 => MR_int_2_26_port, A2 => net134923, ZN => 
                           net60477);
   U665 : NAND2_X1 port map( A1 => n279, A2 => net60477, ZN => MR_int_3_22_port
                           );
   U666 : NAND2_X1 port map( A1 => net61774, A2 => net134969, ZN => n332);
   U667 : NOR2_X1 port map( A1 => net134971, A2 => n385, ZN => n274);
   U668 : NAND2_X1 port map( A1 => ML_int_4_10_port, A2 => net134811, ZN => 
                           n299);
   U669 : NAND2_X1 port map( A1 => ML_int_3_10_port, A2 => net134831, ZN => 
                           n138);
   U670 : NAND2_X1 port map( A1 => ML_int_3_10_port, A2 => net134849, ZN => 
                           n370);
   U671 : NAND2_X1 port map( A1 => n540, A2 => n539, ZN => ML_int_3_10_port);
   U672 : AND2_X1 port map( A1 => n622, A2 => ML_int_4_13_port, ZN => 
                           ML_int_7_13_port);
   U673 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => net134831, ZN => n82)
                           ;
   U674 : NAND2_X1 port map( A1 => n529, A2 => n528, ZN => B(30));
   U675 : NAND2_X1 port map( A1 => n144, A2 => n145, ZN => ML_int_4_26_port);
   U676 : NAND2_X1 port map( A1 => ML_int_3_26_port, A2 => net134831, ZN => 
                           n144);
   U677 : NAND2_X1 port map( A1 => net134861, A2 => n155, ZN => n743);
   U678 : NAND2_X1 port map( A1 => n533, A2 => n534, ZN => n312);
   U679 : AND2_X1 port map( A1 => net60450, A2 => n104, ZN => n99);
   U680 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => net134833, ZN => n81)
                           ;
   U681 : NAND2_X1 port map( A1 => n587, A2 => n586, ZN => ML_int_3_6_port);
   U682 : OAI21_X1 port map( B1 => n219, B2 => net134929, A => n464, ZN => 
                           ML_int_3_23_port);
   U683 : NAND2_X1 port map( A1 => ML_int_2_23_port, A2 => net134929, ZN => 
                           n464);
   U684 : NOR2_X1 port map( A1 => net134831, A2 => n448, ZN => n520);
   U685 : NAND2_X1 port map( A1 => ML_int_3_21_port, A2 => net134849, ZN => 
                           n386);
   U686 : NAND2_X1 port map( A1 => MR_int_4_4_port, A2 => n214, ZN => n212);
   U687 : NAND2_X1 port map( A1 => n345, A2 => net134927, ZN => n465);
   U688 : NAND2_X1 port map( A1 => ML_int_2_9_port, A2 => net134945, ZN => n517
                           );
   U689 : NAND2_X1 port map( A1 => n200, A2 => n505, ZN => n345);
   U690 : NAND2_X1 port map( A1 => MR_int_3_23_port, A2 => net134843, ZN => 
                           n602);
   U691 : NAND2_X1 port map( A1 => MR_int_3_23_port, A2 => n184, ZN => n182);
   U692 : NAND2_X1 port map( A1 => n576, A2 => n577, ZN => B(2));
   U693 : NAND2_X1 port map( A1 => MR_int_5_3_port, A2 => n549, ZN => n576);
   U694 : NAND2_X1 port map( A1 => n314, A2 => n315, ZN => MR_int_5_3_port);
   U695 : NAND2_X1 port map( A1 => ML_int_2_16_port, A2 => net134937, ZN => 
                           n507);
   U696 : NAND2_X1 port map( A1 => ML_int_2_16_port, A2 => net134925, ZN => 
                           n518);
   U697 : NAND2_X1 port map( A1 => n404, A2 => n403, ZN => ML_int_2_16_port);
   U698 : NAND2_X1 port map( A1 => n478, A2 => n479, ZN => MR_int_3_21_port);
   U699 : NAND2_X1 port map( A1 => MR_int_3_21_port, A2 => net134831, ZN => 
                           n338);
   U700 : NAND2_X1 port map( A1 => MR_int_2_20_port, A2 => net134923, ZN => 
                           n591);
   U701 : NAND2_X1 port map( A1 => MR_int_2_20_port, A2 => net134945, ZN => 
                           n566);
   U702 : NAND2_X1 port map( A1 => net61724, A2 => n354, ZN => MR_int_2_20_port
                           );
   U703 : NAND2_X1 port map( A1 => ML_int_2_10_port, A2 => net134927, ZN => 
                           n539);
   U704 : NAND2_X1 port map( A1 => ML_int_2_10_port, A2 => net134947, ZN => 
                           n553);
   U705 : NAND2_X1 port map( A1 => ML_int_2_11_port, A2 => net134925, ZN => 
                           n537);
   U706 : NAND2_X1 port map( A1 => ML_int_2_11_port, A2 => net134941, ZN => 
                           n142);
   U707 : NAND2_X1 port map( A1 => MR_int_4_2_port, A2 => net134809, ZN => n588
                           );
   U708 : NAND2_X1 port map( A1 => n153, A2 => n154, ZN => MR_int_2_2_port);
   U709 : NAND2_X1 port map( A1 => MR_int_1_4_port, A2 => net134879, ZN => n153
                           );
   U710 : NAND2_X1 port map( A1 => n386, A2 => n387, ZN => ML_int_4_29_port);
   U711 : NAND2_X1 port map( A1 => n390, A2 => n389, ZN => ML_int_3_29_port);
   U712 : NAND2_X1 port map( A1 => MR_int_2_29_port, A2 => net134927, ZN => 
                           n147);
   U713 : NAND2_X1 port map( A1 => n445, A2 => n444, ZN => MR_int_3_23_port);
   U714 : NAND2_X1 port map( A1 => MR_int_2_23_port, A2 => net134933, ZN => 
                           n445);
   U715 : NAND2_X1 port map( A1 => MR_int_3_9_port, A2 => n745, ZN => n744);
   U716 : AND2_X1 port map( A1 => net134833, A2 => net134811, ZN => n745);
   U717 : NAND2_X1 port map( A1 => n318, A2 => n319, ZN => B(28));
   U718 : AND2_X1 port map( A1 => net141573, A2 => net134837, ZN => n309);
   U719 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => net134843, ZN => n416
                           );
   U720 : NAND2_X1 port map( A1 => MR_int_1_6_port, A2 => net134899, ZN => n380
                           );
   U721 : NAND2_X1 port map( A1 => n380, A2 => n381, ZN => MR_int_2_6_port);
   U722 : NAND2_X1 port map( A1 => n730, A2 => n175, ZN => n449);
   U723 : AND2_X1 port map( A1 => MR_int_3_24_port, A2 => net134843, ZN => 
                           MR_int_4_24_port);
   U724 : NAND2_X1 port map( A1 => n730, A2 => net134837, ZN => n628);
   U725 : AND2_X1 port map( A1 => net134861, A2 => n155, ZN => MR_int_4_30_port
                           );
   U726 : NOR2_X1 port map( A1 => net134929, A2 => n751, ZN => n155);
   U727 : INV_X1 port map( A => MR_int_2_30_port, ZN => n751);
   U728 : AND2_X1 port map( A1 => n352, A2 => n353, ZN => n219);
   U729 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => ML_int_2_19_port);
   U730 : NAND2_X1 port map( A1 => ML_int_1_19_port, A2 => net135859, ZN => 
                           n352);
   U731 : NAND2_X1 port map( A1 => MR_int_2_11_port, A2 => net134951, ZN => 
                           n554);
   U733 : NAND2_X1 port map( A1 => MR_int_3_7_port, A2 => net134851, ZN => n192
                           );
   U735 : NAND2_X1 port map( A1 => n147, A2 => n148, ZN => MR_int_3_25_port);
   U736 : NAND2_X1 port map( A1 => MR_int_2_27_port, A2 => net134927, ZN => 
                           n444);
   U737 : NAND2_X1 port map( A1 => MR_int_4_3_port, A2 => net134809, ZN => n314
                           );
   U738 : NAND2_X1 port map( A1 => n554, A2 => n555, ZN => MR_int_3_11_port);
   U739 : NAND2_X1 port map( A1 => n511, A2 => n510, ZN => ML_int_3_21_port);
   U740 : NAND2_X1 port map( A1 => n459, A2 => n458, ZN => ML_int_2_21_port);
   U741 : NAND2_X1 port map( A1 => n725, A2 => net134969, ZN => n448);
   U742 : NAND2_X1 port map( A1 => MR_int_3_27_port, A2 => net134831, ZN => 
                           n605);
   U743 : NAND2_X1 port map( A1 => net61842, A2 => n604, ZN => n223);
   U744 : NAND2_X1 port map( A1 => n395, A2 => n396, ZN => ML_int_4_13_port);
   U745 : AND2_X1 port map( A1 => n355, A2 => n356, ZN => n395);
   U746 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => net134845, ZN => n396
                           );
   U747 : NAND2_X1 port map( A1 => n300, A2 => n301, ZN => ML_int_3_5_port);
   U748 : NAND2_X1 port map( A1 => ML_int_2_1_port, A2 => net134943, ZN => n301
                           );
   U749 : NAND2_X1 port map( A1 => net61783, A2 => net61782, ZN => 
                           ML_int_2_20_port);
   U750 : NAND2_X1 port map( A1 => n556, A2 => n557, ZN => MR_int_3_9_port);
   U751 : AND2_X1 port map( A1 => net60450, A2 => n104, ZN => n286);
   U752 : OR2_X1 port map( A1 => n267, A2 => net135875, ZN => n500);
   U753 : NAND2_X1 port map( A1 => MR_int_7_30_port, A2 => net135876, ZN => 
                           n528);
   U754 : NAND2_X1 port map( A1 => MR_int_7_20_port, A2 => net135875, ZN => 
                           n442);
   U755 : NAND2_X1 port map( A1 => MR_int_7_24_port, A2 => net135875, ZN => 
                           n526);
   U756 : NAND2_X1 port map( A1 => n425, A2 => n426, ZN => ML_int_4_19_port);
   U757 : NAND2_X1 port map( A1 => ML_int_3_19_port, A2 => net134851, ZN => 
                           n429);
   U758 : NAND2_X1 port map( A1 => n135, A2 => n136, ZN => MR_int_3_1_port);
   U759 : NAND2_X1 port map( A1 => MR_int_1_5_port, A2 => net134895, ZN => n333
                           );
   U760 : NAND2_X1 port map( A1 => MR_int_4_20_port, A2 => n201, ZN => n213);
   U761 : NAND2_X1 port map( A1 => n522, A2 => n523, ZN => MR_int_4_20_port);
   U762 : NAND2_X1 port map( A1 => n522, A2 => n523, ZN => n156);
   U763 : NAND2_X1 port map( A1 => MR_int_3_20_port, A2 => net134839, ZN => 
                           n522);
   U764 : NAND2_X1 port map( A1 => n551, A2 => n550, ZN => ML_int_4_14_port);
   U765 : NAND2_X1 port map( A1 => n494, A2 => net61053, ZN => ML_int_4_30_port
                           );
   U766 : NAND2_X1 port map( A1 => MR_int_1_16_port, A2 => net134895, ZN => 
                           n542);
   U767 : NAND2_X1 port map( A1 => MR_int_1_16_port, A2 => net134879, ZN => 
                           n283);
   U769 : NAND2_X1 port map( A1 => n542, A2 => net60763, ZN => MR_int_2_16_port
                           );
   U770 : NAND2_X1 port map( A1 => MR_int_2_16_port, A2 => net134923, ZN => 
                           n308);
   U771 : NAND2_X1 port map( A1 => MR_int_2_16_port, A2 => net134949, ZN => 
                           n590);
   U772 : NAND2_X1 port map( A1 => n535, A2 => n536, ZN => MR_int_3_18_port);
   U773 : NAND2_X1 port map( A1 => net61353, A2 => net134947, ZN => n535);
   U774 : NAND2_X1 port map( A1 => n398, A2 => n397, ZN => ML_int_2_10_port);
   U775 : NOR2_X1 port map( A1 => net61363, A2 => net61364, ZN => n100);
   U776 : NOR2_X1 port map( A1 => net61363, A2 => net61364, ZN => n284);
   U778 : NAND2_X1 port map( A1 => n597, A2 => n598, ZN => MR_int_2_29_port);
   U779 : NAND2_X1 port map( A1 => MR_int_1_30_port, A2 => net141464, ZN => 
                           n570);
   U780 : AND2_X1 port map( A1 => net134901, A2 => MR_int_1_30_port, ZN => 
                           MR_int_2_30_port);
   U781 : NAND2_X1 port map( A1 => n97, A2 => net135876, ZN => n91);
   U782 : NAND2_X1 port map( A1 => MR_int_2_1_port, A2 => net134951, ZN => n136
                           );
   U783 : NAND2_X1 port map( A1 => MR_int_4_18_port, A2 => net134969, ZN => 
                           n589);
   U784 : NAND2_X1 port map( A1 => n563, A2 => n562, ZN => MR_int_2_26_port);
   U785 : NAND2_X1 port map( A1 => n527, A2 => n526, ZN => B(24));
   U786 : NAND2_X1 port map( A1 => ML_int_1_14_port, A2 => net134879, ZN => 
                           n508);
   U787 : NAND2_X1 port map( A1 => ML_int_1_14_port, A2 => net134889, ZN => 
                           n404);
   U788 : NAND2_X1 port map( A1 => MR_int_1_25_port, A2 => net134891, ZN => 
                           n543);
   U789 : NAND2_X1 port map( A1 => MR_int_2_9_port, A2 => net134939, ZN => n556
                           );
   U790 : NAND2_X1 port map( A1 => net61046, A2 => n495, ZN => B(22));
   U791 : NOR3_X1 port map( A1 => net134969, A2 => SHMAG_5_port, A3 => n580, ZN
                           => MR_int_7_22_port);
   U792 : NAND2_X1 port map( A1 => MR_int_1_20_port, A2 => net134901, ZN => 
                           net61724);
   U793 : NAND4_X1 port map( A1 => n101, A2 => n98, A3 => n99, A4 => n100, ZN 
                           => n97);
   U794 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => B(10));
   U795 : AOI22_X1 port map( A1 => MR_int_4_11_port, A2 => n383, B1 => n520, B2
                           => n261, ZN => n584);
   U796 : NAND2_X1 port map( A1 => ML_int_7_28_port, A2 => net134977, ZN => 
                           n318);
   U797 : NAND2_X1 port map( A1 => ML_int_7_1_port, A2 => net134977, ZN => n611
                           );
   U798 : NAND2_X1 port map( A1 => ML_int_7_2_port, A2 => net134977, ZN => n577
                           );
   U799 : NAND2_X1 port map( A1 => ML_int_7_6_port, A2 => net134977, ZN => n461
                           );
   U800 : NAND2_X1 port map( A1 => ML_int_7_0_port, A2 => net134977, ZN => n502
                           );
   U801 : NAND2_X1 port map( A1 => ML_int_7_3_port, A2 => net134977, ZN => n583
                           );
   U802 : NAND2_X1 port map( A1 => ML_int_7_14_port, A2 => net134977, ZN => 
                           n569);
   U803 : NAND2_X1 port map( A1 => ML_int_7_10_port, A2 => net134977, ZN => 
                           n585);
   U804 : NAND2_X1 port map( A1 => ML_int_7_7_port, A2 => net134977, ZN => n477
                           );
   U805 : NAND2_X1 port map( A1 => n560, A2 => n561, ZN => MR_int_2_22_port);
   U806 : NAND2_X1 port map( A1 => MR_int_2_22_port, A2 => net134925, ZN => 
                           n536);
   U807 : NAND2_X1 port map( A1 => MR_int_2_22_port, A2 => net134947, ZN => 
                           n279);
   U808 : NAND2_X1 port map( A1 => MR_int_2_15_port, A2 => net134943, ZN => 
                           n346);
   U809 : NAND2_X1 port map( A1 => MR_int_2_15_port, A2 => net134923, ZN => 
                           n555);
   U810 : NAND2_X1 port map( A1 => n581, A2 => net60604, ZN => MR_int_2_15_port
                           );
   U811 : NAND2_X1 port map( A1 => MR_int_2_5_port, A2 => net134929, ZN => n135
                           );
   U812 : NAND2_X1 port map( A1 => n333, A2 => n334, ZN => MR_int_2_5_port);
   U813 : NAND2_X1 port map( A1 => n726, A2 => net134843, ZN => n197);
   U814 : NAND2_X1 port map( A1 => n236, A2 => net134831, ZN => net61842);
   U815 : NAND2_X1 port map( A1 => n178, A2 => n255, ZN => B(7));
   U816 : NAND2_X1 port map( A1 => MR_int_1_29_port, A2 => net134899, ZN => 
                           n597);
   U817 : NAND2_X1 port map( A1 => n347, A2 => n346, ZN => MR_int_3_15_port);
   U818 : NAND2_X1 port map( A1 => MR_int_2_24_port, A2 => net134941, ZN => 
                           n485);
   U819 : NAND2_X1 port map( A1 => MR_int_2_24_port, A2 => net134925, ZN => 
                           n567);
   U820 : NAND2_X1 port map( A1 => n332, A2 => n331, ZN => n181);
   U821 : NAND2_X1 port map( A1 => MR_int_4_6_port, A2 => net134809, ZN => n331
                           );
   U822 : NAND2_X1 port map( A1 => MR_int_2_14_port, A2 => net134947, ZN => 
                           net60589);
   U823 : NAND2_X1 port map( A1 => MR_int_2_14_port, A2 => net134923, ZN => 
                           net61331);
   U824 : NAND2_X1 port map( A1 => n283, A2 => n282, ZN => MR_int_2_14_port);
   U825 : NAND2_X1 port map( A1 => n599, A2 => n600, ZN => MR_int_2_24_port);
   U826 : NAND2_X1 port map( A1 => MR_int_1_26_port, A2 => net134895, ZN => 
                           n562);
   U827 : AND2_X1 port map( A1 => n578, A2 => n665, ZN => n224);
   U828 : NAND2_X1 port map( A1 => MR_int_2_25_port, A2 => net134935, ZN => 
                           n148);
   U829 : NAND2_X1 port map( A1 => MR_int_2_25_port, A2 => net134927, ZN => 
                           n479);
   U830 : NAND2_X1 port map( A1 => n543, A2 => n544, ZN => MR_int_2_25_port);
   U831 : NAND2_X1 port map( A1 => MR_int_3_9_port, A2 => net134843, ZN => n467
                           );
   U832 : NAND2_X1 port map( A1 => ML_int_3_18_port, A2 => net134833, ZN => 
                           n369);
   U833 : NAND2_X1 port map( A1 => n521, A2 => net60893, ZN => ML_int_3_18_port
                           );
   U834 : NAND2_X1 port map( A1 => MR_int_1_10_port, A2 => net134875, ZN => 
                           n498);
   U835 : NAND2_X1 port map( A1 => MR_int_1_18_port, A2 => net141528, ZN => 
                           net60763);
   U836 : NAND2_X1 port map( A1 => MR_int_1_8_port, A2 => net141464, ZN => n381
                           );
   U837 : NAND2_X1 port map( A1 => n186, A2 => net134875, ZN => n354);
   U838 : NAND2_X1 port map( A1 => ML_int_1_4_port, A2 => net135858, ZN => 
                           net60869);
   U839 : NAND2_X1 port map( A1 => ML_int_1_8_port, A2 => net135858, ZN => n334
                           );
   U840 : NAND2_X1 port map( A1 => ML_int_1_22_port, A2 => net135858, ZN => 
                           n311);
   U841 : NAND2_X1 port map( A1 => ML_int_1_2_port, A2 => net141528, ZN => n195
                           );
   U842 : NAND2_X1 port map( A1 => ML_int_1_18_port, A2 => net135858, ZN => 
                           n326);
   U843 : NOR2_X1 port map( A1 => net60750, A2 => net60751, ZN => n101);
   U844 : NOR2_X1 port map( A1 => net60750, A2 => net60751, ZN => n285);
   U845 : NAND2_X1 port map( A1 => MR_int_2_21_port, A2 => net134927, ZN => 
                           n565);
   U846 : AND2_X1 port map( A1 => n574, A2 => n575, ZN => n541);
   U847 : NAND2_X1 port map( A1 => n660, A2 => n575, ZN => MR_int_4_18_port);
   U848 : NAND2_X1 port map( A1 => MR_int_7_22_port, A2 => net135876, ZN => 
                           net61046);
   U849 : NAND2_X1 port map( A1 => n564, A2 => n565, ZN => MR_int_3_17_port);
   U850 : NAND2_X1 port map( A1 => n264, A2 => net134933, ZN => net61039);
   U851 : NAND2_X1 port map( A1 => n496, A2 => net61039, ZN => ML_int_3_17_port
                           );
   U852 : NAND2_X1 port map( A1 => ML_int_4_17_port, A2 => net134821, ZN => 
                           n360);
   U853 : NAND2_X1 port map( A1 => n351, A2 => n350, ZN => ML_int_2_11_port);
   U854 : NAND2_X1 port map( A1 => ML_int_1_9_port, A2 => net134889, ZN => n351
                           );
   U855 : NAND2_X1 port map( A1 => n514, A2 => n515, ZN => B(23));
   U856 : NAND2_X1 port map( A1 => n571, A2 => n570, ZN => n623);
   U857 : AND2_X1 port map( A1 => n570, A2 => n571, ZN => n215);
   U858 : NAND2_X1 port map( A1 => n336, A2 => n335, ZN => B(25));
   U859 : NOR2_X1 port map( A1 => net65464, A2 => net65465, ZN => n98);
   U860 : NOR2_X1 port map( A1 => net65464, A2 => net65465, ZN => n270);
   U861 : NAND2_X1 port map( A1 => n411, A2 => n412, ZN => n272);
   U862 : NAND2_X1 port map( A1 => MR_int_3_17_port, A2 => net134839, ZN => 
                           n579);
   U863 : NAND2_X1 port map( A1 => MR_int_3_15_port, A2 => net134851, ZN => 
                           n422);
   U864 : NAND2_X1 port map( A1 => MR_int_3_15_port, A2 => net134831, ZN => 
                           n193);
   U865 : NAND2_X1 port map( A1 => MR_int_2_19_port, A2 => net134949, ZN => 
                           n546);
   U866 : NAND2_X1 port map( A1 => MR_int_2_19_port, A2 => net134925, ZN => 
                           n347);
   U867 : NAND2_X1 port map( A1 => MR_int_3_25_port, A2 => net134833, ZN => 
                           n243);
   U868 : AND2_X1 port map( A1 => MR_int_3_25_port, A2 => net134839, ZN => 
                           MR_int_4_25_port);
   U869 : NAND2_X1 port map( A1 => MR_int_3_25_port, A2 => net134833, ZN => 
                           n578);
   U870 : NAND2_X1 port map( A1 => MR_int_1_24_port, A2 => net141528, ZN => 
                           n560);
   U871 : NAND2_X1 port map( A1 => n482, A2 => n483, ZN => ML_int_2_12_port);
   U872 : NAND2_X1 port map( A1 => ML_int_1_12_port, A2 => net134879, ZN => 
                           n482);
   U873 : NAND2_X1 port map( A1 => n321, A2 => n320, ZN => n251);
   U874 : NAND2_X1 port map( A1 => ML_int_2_8_port, A2 => net134937, ZN => n321
                           );
   U875 : NAND2_X1 port map( A1 => MR_int_4_19_port, A2 => net134821, ZN => 
                           n315);
   U876 : NAND2_X1 port map( A1 => n605, A2 => n604, ZN => MR_int_4_19_port);
   U877 : NAND2_X1 port map( A1 => MR_int_3_19_port, A2 => net134839, ZN => 
                           n604);
   U878 : NAND2_X1 port map( A1 => n545, A2 => n546, ZN => MR_int_3_19_port);
   U879 : NAND2_X1 port map( A1 => n558, A2 => n559, ZN => B(5));
   U880 : NAND4_X1 port map( A1 => n285, A2 => n286, A3 => n284, A4 => n270, ZN
                           => net60578);
   U881 : NAND2_X1 port map( A1 => ML_int_3_19_port, A2 => net134831, ZN => 
                           n425);
   U882 : NAND2_X1 port map( A1 => ML_int_2_19_port, A2 => net134925, ZN => 
                           n503);
   U883 : AND2_X1 port map( A1 => MR_int_3_26_port, A2 => net134839, ZN => n229
                           );
   U884 : NAND2_X1 port map( A1 => net134855, A2 => MR_int_3_26_port, ZN => 
                           n385);
   U885 : NAND2_X1 port map( A1 => MR_int_3_26_port, A2 => net134833, ZN => 
                           n574);
   U886 : NAND2_X1 port map( A1 => n732, A2 => net134883, ZN => n571);
   U887 : AND2_X1 port map( A1 => net135715, A2 => n90, ZN => n173);
   U888 : NAND2_X1 port map( A1 => MR_int_1_28_port, A2 => net141528, ZN => 
                           n563);
   U889 : NAND2_X1 port map( A1 => net135715, A2 => n90, ZN => 
                           temp_int_SH_4_port);
   U890 : AND2_X1 port map( A1 => n695, A2 => A(0), ZN => ML_int_1_0_port);
   U891 : NOR2_X1 port map( A1 => n749, A2 => net141178, ZN => MR_int_1_31_port
                           );
   U892 : NAND2_X1 port map( A1 => ML_int_2_21_port, A2 => net134949, ZN => 
                           n487);
   U893 : NAND2_X1 port map( A1 => MR_int_1_26_port, A2 => net135859, ZN => 
                           n600);
   U894 : NAND2_X1 port map( A1 => ML_int_1_16_port, A2 => net134875, ZN => 
                           n403);
   U895 : NAND2_X1 port map( A1 => ML_int_1_23_port, A2 => net134875, ZN => 
                           n121);
   U896 : NAND2_X1 port map( A1 => ML_int_1_6_port, A2 => net135858, ZN => n393
                           );
   U897 : NAND2_X1 port map( A1 => ML_int_1_11_port, A2 => net135858, ZN => 
                           n350);
   U898 : NAND2_X1 port map( A1 => ML_int_1_20_port, A2 => net135858, ZN => 
                           net61782);
   U899 : NAND2_X1 port map( A1 => ML_int_1_10_port, A2 => net135859, ZN => 
                           n397);
   U900 : NAND2_X1 port map( A1 => MR_int_1_21_port, A2 => net134875, ZN => 
                           n596);
   U901 : NAND2_X1 port map( A1 => MR_int_1_27_port, A2 => net141528, ZN => 
                           n544);
   U902 : NAND2_X1 port map( A1 => n601, A2 => net135859, ZN => n609);
   U903 : NAND2_X1 port map( A1 => ML_int_1_21_port, A2 => net135858, ZN => 
                           n458);
   U904 : INV_X2 port map( A => net134859, ZN => net134831);
   U905 : AND2_X4 port map( A1 => net135715, A2 => n92, ZN => SHMAG_5_port);
   U906 : INV_X1 port map( A => net134825, ZN => net134813);
   U907 : INV_X1 port map( A => temp_int_SH_4_port, ZN => net134815);
   U908 : INV_X1 port map( A => temp_int_SH_4_port, ZN => net134819);
   U909 : INV_X1 port map( A => temp_int_SH_4_port, ZN => net134821);
   U910 : INV_X1 port map( A => temp_int_SH_4_port, ZN => net134825);
   U911 : INV_X1 port map( A => temp_int_SH_4_port, ZN => net134827);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity COMPARATOR_M32 is

   port( A, B : in std_logic_vector (31 downto 0);  sel : in std_logic_vector 
         (1 downto 0);  OUTPUT : out std_logic_vector (31 downto 0));

end COMPARATOR_M32;

architecture SYN_BEHAVIORAL of COMPARATOR_M32 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component COMPARATOR_M32_DW01_cmp6_1
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, OUTPUT_0_port, N12, N15, N16, n1, n5, n6, n8, n9, 
      n_1024, n_1025, n_1026 : std_logic;

begin
   OUTPUT <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      OUTPUT_0_port );
   
   X_Logic0_port <= '0';
   n1 <= '0';
   U8 : XOR2_X1 port map( A => n8, B => N12, Z => n6);
   r61 : COMPARATOR_M32_DW01_cmp6_1 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), TC => n1, LT => n_1024, GT => 
                           n_1025, EQ => N12, LE => N16, GE => N15, NE => 
                           n_1026);
   U2 : INV_X1 port map( A => sel(1), ZN => n9);
   U4 : AOI22_X1 port map( A1 => N15, A2 => n8, B1 => N16, B2 => sel(0), ZN => 
                           n5);
   U5 : INV_X1 port map( A => sel(0), ZN => n8);
   U6 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => sel(1), B2 => n6, ZN => 
                           OUTPUT_0_port);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity P4ADDER_n_bit32 is

   port( A, B : in std_logic_vector (31 downto 0);  cin0 : in std_logic;  S : 
         out std_logic_vector (31 downto 0));

end P4ADDER_n_bit32;

architecture SYN_STRUCTURAL of P4ADDER_n_bit32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CSA
      port( A, B : in std_logic_vector (31 downto 0);  c : in std_logic_vector 
            (7 downto 0);  s : out std_logic_vector (31 downto 0));
   end component;
   
   component Cg
      port( A, B : in std_logic_vector (31 downto 0);  cin0 : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carries_7_port, carries_6_port, carries_5_port, carries_4_port, 
      carries_3_port, carries_2_port, carries_1_port, BS_31_port, BS_30_port, 
      BS_29_port, BS_28_port, BS_27_port, BS_26_port, BS_25_port, BS_24_port, 
      BS_23_port, BS_22_port, BS_21_port, BS_20_port, BS_19_port, BS_18_port, 
      BS_17_port, BS_16_port, BS_15_port, BS_14_port, BS_13_port, BS_12_port, 
      BS_11_port, BS_10_port, BS_9_port, BS_8_port, BS_7_port, BS_6_port, 
      BS_5_port, BS_4_port, BS_3_port, BS_2_port, BS_1_port, n1, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n_1027 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n17, B => B(8), Z => BS_8_port);
   U4 : XOR2_X1 port map( A => n17, B => B(7), Z => BS_7_port);
   U5 : XOR2_X1 port map( A => n17, B => B(6), Z => BS_6_port);
   U6 : XOR2_X1 port map( A => n17, B => B(5), Z => BS_5_port);
   U7 : XOR2_X1 port map( A => n17, B => B(4), Z => BS_4_port);
   U9 : XOR2_X1 port map( A => n17, B => B(31), Z => BS_31_port);
   U10 : XOR2_X1 port map( A => n17, B => B(30), Z => BS_30_port);
   U11 : XOR2_X1 port map( A => n17, B => B(2), Z => BS_2_port);
   U12 : XOR2_X1 port map( A => n17, B => B(29), Z => BS_29_port);
   U13 : XOR2_X1 port map( A => n17, B => B(28), Z => BS_28_port);
   U14 : XOR2_X1 port map( A => n17, B => B(27), Z => BS_27_port);
   U15 : XOR2_X1 port map( A => n17, B => B(26), Z => BS_26_port);
   U16 : XOR2_X1 port map( A => n17, B => B(25), Z => BS_25_port);
   U17 : XOR2_X1 port map( A => n17, B => B(24), Z => BS_24_port);
   U18 : XOR2_X1 port map( A => n17, B => B(23), Z => BS_23_port);
   U19 : XOR2_X1 port map( A => n17, B => B(22), Z => BS_22_port);
   U20 : XOR2_X1 port map( A => n17, B => B(21), Z => BS_21_port);
   U21 : XOR2_X1 port map( A => n17, B => B(20), Z => BS_20_port);
   U22 : XOR2_X1 port map( A => n17, B => B(1), Z => BS_1_port);
   U23 : XOR2_X1 port map( A => n17, B => B(19), Z => BS_19_port);
   U24 : XOR2_X1 port map( A => n17, B => B(18), Z => BS_18_port);
   U25 : XOR2_X1 port map( A => n17, B => B(17), Z => BS_17_port);
   U26 : XOR2_X1 port map( A => n17, B => B(16), Z => BS_16_port);
   U27 : XOR2_X1 port map( A => n17, B => B(15), Z => BS_15_port);
   U28 : XOR2_X1 port map( A => n17, B => B(14), Z => BS_14_port);
   U29 : XOR2_X1 port map( A => n17, B => B(13), Z => BS_13_port);
   U30 : XOR2_X1 port map( A => n17, B => B(12), Z => BS_12_port);
   U31 : XOR2_X1 port map( A => n17, B => B(11), Z => BS_11_port);
   U32 : XOR2_X1 port map( A => n17, B => B(10), Z => BS_10_port);
   CG1 : Cg port map( A(31) => A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => BS_31_port, B(30) => BS_30_port, B(29) => 
                           BS_29_port, B(28) => BS_28_port, B(27) => BS_27_port
                           , B(26) => BS_26_port, B(25) => BS_25_port, B(24) =>
                           BS_24_port, B(23) => BS_23_port, B(22) => BS_22_port
                           , B(21) => BS_21_port, B(20) => BS_20_port, B(19) =>
                           BS_19_port, B(18) => BS_18_port, B(17) => BS_17_port
                           , B(16) => BS_16_port, B(15) => BS_15_port, B(14) =>
                           BS_14_port, B(13) => BS_13_port, B(12) => BS_12_port
                           , B(11) => BS_11_port, B(10) => BS_10_port, B(9) => 
                           BS_9_port, B(8) => BS_8_port, B(7) => BS_7_port, 
                           B(6) => BS_6_port, B(5) => BS_5_port, B(4) => 
                           BS_4_port, B(3) => BS_3_port, B(2) => BS_2_port, 
                           B(1) => BS_1_port, B(0) => n1, cin0 => n17, cout(7) 
                           => n_1027, cout(6) => carries_7_port, cout(5) => 
                           carries_6_port, cout(4) => carries_5_port, cout(3) 
                           => carries_4_port, cout(2) => carries_3_port, 
                           cout(1) => carries_2_port, cout(0) => carries_1_port
                           );
   CSA1 : CSA port map( A(31) => A(31), A(30) => A(30), A(29) => A(29), A(28) 
                           => A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => BS_31_port, B(30) => BS_30_port, B(29) => 
                           BS_29_port, B(28) => BS_28_port, B(27) => BS_27_port
                           , B(26) => BS_26_port, B(25) => BS_25_port, B(24) =>
                           BS_24_port, B(23) => BS_23_port, B(22) => BS_22_port
                           , B(21) => BS_21_port, B(20) => BS_20_port, B(19) =>
                           BS_19_port, B(18) => BS_18_port, B(17) => BS_17_port
                           , B(16) => BS_16_port, B(15) => n15, B(14) => n5, 
                           B(13) => n7, B(12) => BS_12_port, B(11) => n14, 
                           B(10) => BS_10_port, B(9) => n13, B(8) => BS_8_port,
                           B(7) => n6, B(6) => BS_6_port, B(5) => n4, B(4) => 
                           BS_4_port, B(3) => n12, B(2) => BS_2_port, B(1) => 
                           n11, B(0) => n16, c(7) => carries_7_port, c(6) => 
                           carries_6_port, c(5) => carries_5_port, c(4) => 
                           carries_4_port, c(3) => carries_3_port, c(2) => 
                           carries_2_port, c(1) => carries_1_port, c(0) => n17,
                           s(31) => S(31), s(30) => S(30), s(29) => S(29), 
                           s(28) => S(28), s(27) => S(27), s(26) => S(26), 
                           s(25) => S(25), s(24) => S(24), s(23) => S(23), 
                           s(22) => S(22), s(21) => S(21), s(20) => S(20), 
                           s(19) => S(19), s(18) => S(18), s(17) => S(17), 
                           s(16) => S(16), s(15) => S(15), s(14) => S(14), 
                           s(13) => S(13), s(12) => S(12), s(11) => S(11), 
                           s(10) => S(10), s(9) => S(9), s(8) => S(8), s(7) => 
                           S(7), s(6) => S(6), s(5) => S(5), s(4) => S(4), s(3)
                           => S(3), s(2) => S(2), s(1) => S(1), s(0) => S(0));
   U1 : BUF_X4 port map( A => cin0, Z => n17);
   U2 : CLKBUF_X1 port map( A => BS_5_port, Z => n4);
   U8 : XNOR2_X1 port map( A => n8, B => B(9), ZN => BS_9_port);
   U33 : XNOR2_X1 port map( A => n8, B => B(0), ZN => n1);
   U34 : XOR2_X1 port map( A => n17, B => B(14), Z => n5);
   U35 : XOR2_X1 port map( A => n17, B => B(7), Z => n6);
   U36 : XOR2_X1 port map( A => n17, B => B(13), Z => n7);
   U37 : OR2_X1 port map( A1 => B(3), A2 => n8, ZN => n9);
   U38 : INV_X1 port map( A => cin0, ZN => n8);
   U39 : NAND2_X1 port map( A1 => B(3), A2 => n8, ZN => n10);
   U40 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => BS_3_port);
   U41 : CLKBUF_X1 port map( A => BS_1_port, Z => n11);
   U42 : CLKBUF_X1 port map( A => BS_3_port, Z => n12);
   U43 : CLKBUF_X1 port map( A => n1, Z => n16);
   U44 : BUF_X1 port map( A => BS_9_port, Z => n13);
   U45 : BUF_X1 port map( A => BS_11_port, Z => n14);
   U46 : BUF_X1 port map( A => BS_15_port, Z => n15);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity SHIFTER_M32_N5 is

   port( A, B : in std_logic_vector (31 downto 0);  LEFT_RIGHT : in std_logic; 
         OUTPUT : out std_logic_vector (31 downto 0));

end SHIFTER_M32_N5;

architecture SYN_BEHAVIORAL of SHIFTER_M32_N5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SHIFTER_M32_N5_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (31 downto 0);  SH_TC : in std_logic;  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_M32_N5_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (31 downto 0);  SH_TC : in std_logic;  B : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31
      , N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, 
      N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60
      , N61, N62, N63, N64, N65, n1, n2_port, n3_port, n4_port, n42_port, 
      n44_port, n49_port, n50_port, n52_port, n53_port, n57_port, n58_port, 
      n59_port, n61_port, n63_port, n64_port, n67, n68, n70, n71, n72, n73, 
      net133051, net133049, net133047, net133045, net133043, net133041, 
      net133037, net133033, net133065, n140, n142, n143, n144, n145, n146, n147
      : std_logic;

begin
   
   n1 <= '1';
   n2_port <= '0';
   n3_port <= '1';
   n4_port <= '0';
   sll_29 : SHIFTER_M32_N5_DW01_ash_0 port map( A(31) => A(31), A(30) => A(30),
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), DATA_TC => n4_port, SH(31) => 
                           B(31), SH(30) => B(30), SH(29) => B(29), SH(28) => 
                           B(28), SH(27) => B(27), SH(26) => B(26), SH(25) => 
                           B(25), SH(24) => B(24), SH(23) => B(23), SH(22) => 
                           B(22), SH(21) => B(21), SH(20) => B(20), SH(19) => 
                           B(19), SH(18) => B(18), SH(17) => B(17), SH(16) => 
                           B(16), SH(15) => B(15), SH(14) => B(14), SH(13) => 
                           B(13), SH(12) => B(12), SH(11) => B(11), SH(10) => 
                           B(10), SH(9) => B(9), SH(8) => B(8), SH(7) => B(7), 
                           SH(6) => B(6), SH(5) => B(5), SH(4) => B(4), SH(3) 
                           => B(3), SH(2) => B(2), SH(1) => B(1), SH(0) => B(0)
                           , SH_TC => n1, B(31) => N65, B(30) => N64, B(29) => 
                           N63, B(28) => N62, B(27) => N61, B(26) => N60, B(25)
                           => N59, B(24) => N58, B(23) => N57, B(22) => N56, 
                           B(21) => N55, B(20) => N54, B(19) => N53, B(18) => 
                           N52, B(17) => N51, B(16) => N50, B(15) => N49, B(14)
                           => N48, B(13) => N47, B(12) => N46, B(11) => N45, 
                           B(10) => N44, B(9) => N43, B(8) => N42, B(7) => N41,
                           B(6) => N40, B(5) => N39, B(4) => N38, B(3) => N37, 
                           B(2) => N36, B(1) => N35, B(0) => N34);
   srl_27 : SHIFTER_M32_N5_DW_rash_0 port map( A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), DATA_TC => n2_port, SH(31) => 
                           B(31), SH(30) => B(30), SH(29) => B(29), SH(28) => 
                           B(28), SH(27) => B(27), SH(26) => B(26), SH(25) => 
                           B(25), SH(24) => B(24), SH(23) => B(23), SH(22) => 
                           B(22), SH(21) => B(21), SH(20) => B(20), SH(19) => 
                           B(19), SH(18) => B(18), SH(17) => B(17), SH(16) => 
                           B(16), SH(15) => B(15), SH(14) => B(14), SH(13) => 
                           B(13), SH(12) => B(12), SH(11) => B(11), SH(10) => 
                           B(10), SH(9) => B(9), SH(8) => B(8), SH(7) => B(7), 
                           SH(6) => B(6), SH(5) => B(5), SH(4) => B(4), SH(3) 
                           => B(3), SH(2) => B(2), SH(1) => B(1), SH(0) => B(0)
                           , SH_TC => n3_port, B(31) => N33, B(30) => N32, 
                           B(29) => N31, B(28) => N30, B(27) => N29, B(26) => 
                           N28, B(25) => N27, B(24) => N26, B(23) => N25, B(22)
                           => N24, B(21) => N23, B(20) => N22, B(19) => N21, 
                           B(18) => N20, B(17) => N19, B(16) => N18, B(15) => 
                           N17, B(14) => N16, B(13) => N15, B(12) => N14, B(11)
                           => N13, B(10) => N12, B(9) => N11, B(8) => N10, B(7)
                           => N9, B(6) => N8, B(5) => N7, B(4) => N6, B(3) => 
                           N5, B(2) => N4, B(1) => N3, B(0) => N2);
   U1 : MUX2_X1 port map( A => N47, B => N15, S => net133033, Z => OUTPUT(13));
   U2 : INV_X1 port map( A => N10, ZN => n140);
   U7 : NAND2_X1 port map( A1 => n142, A2 => n143, ZN => OUTPUT(8));
   U8 : OR2_X1 port map( A1 => n144, A2 => n140, ZN => n142);
   U9 : NAND2_X1 port map( A1 => net133043, A2 => N42, ZN => n143);
   U10 : MUX2_X1 port map( A => N55, B => N23, S => net133033, Z => OUTPUT(21))
                           ;
   U11 : MUX2_X1 port map( A => N38, B => N6, S => net133033, Z => OUTPUT(4));
   U12 : MUX2_X1 port map( A => N5, B => N37, S => LEFT_RIGHT, Z => OUTPUT(3));
   U13 : MUX2_X1 port map( A => N27, B => N59, S => LEFT_RIGHT, Z => OUTPUT(25)
                           );
   U14 : MUX2_X1 port map( A => N29, B => N61, S => LEFT_RIGHT, Z => OUTPUT(27)
                           );
   U15 : MUX2_X1 port map( A => N7, B => N39, S => LEFT_RIGHT, Z => OUTPUT(5));
   U16 : MUX2_X1 port map( A => N8, B => N40, S => LEFT_RIGHT, Z => OUTPUT(6));
   U17 : MUX2_X1 port map( A => N28, B => N60, S => LEFT_RIGHT, Z => OUTPUT(26)
                           );
   U18 : MUX2_X1 port map( A => N18, B => N50, S => LEFT_RIGHT, Z => OUTPUT(16)
                           );
   U19 : MUX2_X1 port map( A => N19, B => N51, S => LEFT_RIGHT, Z => OUTPUT(17)
                           );
   U20 : MUX2_X1 port map( A => N4, B => N36, S => LEFT_RIGHT, Z => OUTPUT(2));
   U21 : MUX2_X1 port map( A => N3, B => N35, S => LEFT_RIGHT, Z => OUTPUT(1));
   U22 : BUF_X1 port map( A => n146, Z => n144);
   U23 : AOI22_X1 port map( A1 => N33, A2 => net133033, B1 => N65, B2 => n144, 
                           ZN => n49_port);
   U24 : BUF_X1 port map( A => LEFT_RIGHT, Z => n146);
   U25 : BUF_X1 port map( A => n146, Z => net133041);
   U26 : BUF_X1 port map( A => n146, Z => net133037);
   U27 : BUF_X1 port map( A => n147, Z => n145);
   U28 : INV_X1 port map( A => n145, ZN => net133033);
   U29 : BUF_X1 port map( A => LEFT_RIGHT, Z => n147);
   U30 : BUF_X1 port map( A => n147, Z => net133049);
   U31 : BUF_X1 port map( A => n147, Z => net133051);
   U32 : BUF_X1 port map( A => LEFT_RIGHT, Z => net133065);
   U33 : BUF_X1 port map( A => net133065, Z => net133045);
   U34 : BUF_X1 port map( A => net133065, Z => net133047);
   U35 : BUF_X1 port map( A => net133065, Z => net133043);
   U36 : AOI22_X1 port map( A1 => N25, A2 => net133033, B1 => N57, B2 => 
                           net133045, ZN => n58_port);
   U37 : INV_X1 port map( A => n44_port, ZN => OUTPUT(7));
   U38 : INV_X1 port map( A => n49_port, ZN => OUTPUT(31));
   U39 : INV_X1 port map( A => n58_port, ZN => OUTPUT(23));
   U40 : INV_X1 port map( A => n68, ZN => OUTPUT(14));
   U41 : INV_X1 port map( A => n63_port, ZN => OUTPUT(19));
   U42 : AOI22_X1 port map( A1 => N24, A2 => net133033, B1 => N56, B2 => 
                           net133045, ZN => n59_port);
   U43 : AOI22_X1 port map( A1 => N30, A2 => net133033, B1 => N62, B2 => 
                           net133041, ZN => n53_port);
   U44 : AOI22_X1 port map( A1 => N16, A2 => net133033, B1 => N48, B2 => 
                           net133049, ZN => n68);
   U45 : AOI22_X1 port map( A1 => N22, A2 => net133033, B1 => N54, B2 => 
                           net133045, ZN => n61_port);
   U46 : AOI22_X1 port map( A1 => N20, A2 => net133033, B1 => N52, B2 => 
                           net133047, ZN => n64_port);
   U47 : AOI22_X1 port map( A1 => N21, A2 => net133033, B1 => N53, B2 => 
                           net133047, ZN => n63_port);
   U48 : INV_X1 port map( A => n61_port, ZN => OUTPUT(20));
   U49 : AOI22_X1 port map( A1 => N13, A2 => net133033, B1 => N45, B2 => 
                           net133051, ZN => n71);
   U50 : INV_X1 port map( A => n52_port, ZN => OUTPUT(29));
   U51 : AOI22_X1 port map( A1 => N14, A2 => net133033, B1 => N46, B2 => 
                           net133051, ZN => n70);
   U52 : AOI22_X1 port map( A1 => N17, A2 => net133033, B1 => N49, B2 => 
                           net133049, ZN => n67);
   U53 : INV_X1 port map( A => n67, ZN => OUTPUT(15));
   U54 : INV_X1 port map( A => n42_port, ZN => OUTPUT(9));
   U55 : AOI22_X1 port map( A1 => N11, A2 => net133033, B1 => N43, B2 => 
                           net133037, ZN => n42_port);
   U56 : INV_X1 port map( A => n59_port, ZN => OUTPUT(22));
   U57 : AOI22_X1 port map( A1 => N32, A2 => net133033, B1 => N64, B2 => 
                           net133041, ZN => n50_port);
   U58 : INV_X1 port map( A => n72, ZN => OUTPUT(10));
   U59 : INV_X1 port map( A => n57_port, ZN => OUTPUT(24));
   U60 : INV_X1 port map( A => n71, ZN => OUTPUT(11));
   U61 : INV_X1 port map( A => n64_port, ZN => OUTPUT(18));
   U62 : INV_X1 port map( A => n50_port, ZN => OUTPUT(30));
   U63 : AOI22_X1 port map( A1 => N26, A2 => net133033, B1 => N58, B2 => 
                           net133043, ZN => n57_port);
   U64 : AOI22_X1 port map( A1 => N12, A2 => net133033, B1 => N44, B2 => 
                           net133051, ZN => n72);
   U65 : INV_X1 port map( A => n70, ZN => OUTPUT(12));
   U66 : AOI22_X1 port map( A1 => N2, A2 => net133033, B1 => N34, B2 => 
                           net133051, ZN => n73);
   U67 : AOI22_X1 port map( A1 => N9, A2 => net133033, B1 => N41, B2 => 
                           net133037, ZN => n44_port);
   U68 : INV_X1 port map( A => n73, ZN => OUTPUT(0));
   U69 : INV_X1 port map( A => n53_port, ZN => OUTPUT(28));
   U70 : AOI22_X1 port map( A1 => N31, A2 => net133033, B1 => N63, B2 => 
                           net133041, ZN => n52_port);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Adder_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end Adder_DW01_add_0;

architecture SYN_rpl of Adder_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, n_1029 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           n_1029, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_6 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_6;

architecture SYN_behavioral of reg_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94
      , n95, n96, n97, n98, n99, n102, net134801, net134799, net134797, 
      net134807, net134805, net134803, n35, n34, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204 : std_logic;

begin
   
   temp_reg_27_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_24_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_22_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_18_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_11_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_8_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n102, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_2_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_0_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(0), QN => 
                           n36);
   temp_reg_23_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_25_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_3_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_13_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_1_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_9_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_20_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_12_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_28_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_31_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_29_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_30_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(30), QN =>
                           n66);
   U3 : BUF_X1 port map( A => n35, Z => net134807);
   U4 : BUF_X1 port map( A => n34, Z => net134801);
   U5 : BUF_X1 port map( A => n35, Z => net134805);
   U6 : BUF_X1 port map( A => n34, Z => net134799);
   U7 : BUF_X1 port map( A => n35, Z => net134803);
   U8 : BUF_X1 port map( A => n34, Z => net134797);
   U9 : OAI22_X1 port map( A1 => n176, A2 => n34, B1 => n35, B2 => n45, ZN => 
                           n89);
   U10 : OAI22_X1 port map( A1 => n202, A2 => n34, B1 => n35, B2 => n42, ZN => 
                           n102);
   U11 : OAI22_X1 port map( A1 => n180, A2 => n34, B1 => n35, B2 => n49, ZN => 
                           n85);
   U12 : OAI22_X1 port map( A1 => n185, A2 => n34, B1 => n35, B2 => n52, ZN => 
                           n82);
   U13 : OAI22_X1 port map( A1 => n190, A2 => n34, B1 => n35, B2 => n63, ZN => 
                           n71);
   U14 : OAI22_X1 port map( A1 => n191, A2 => n34, B1 => n35, B2 => n62, ZN => 
                           n72);
   U15 : OAI22_X1 port map( A1 => n184, A2 => n34, B1 => n35, B2 => n53, ZN => 
                           n81);
   U16 : OAI22_X1 port map( A1 => n188, A2 => n34, B1 => n35, B2 => n57, ZN => 
                           n77);
   U17 : OAI22_X1 port map( A1 => n172, A2 => n34, B1 => n35, B2 => n40, ZN => 
                           n94);
   U18 : INV_X1 port map( A => i(4), ZN => n172);
   U19 : OR2_X1 port map( A1 => reset, A2 => load, ZN => n35);
   U20 : NAND2_X1 port map( A1 => load, A2 => n173, ZN => n34);
   U21 : INV_X1 port map( A => reset, ZN => n173);
   U22 : OAI22_X1 port map( A1 => net134799, A2 => n178, B1 => net134805, B2 =>
                           n51, ZN => n83);
   U23 : INV_X1 port map( A => i(10), ZN => n175);
   U24 : OAI22_X1 port map( A1 => net134801, A2 => n194, B1 => net134807, B2 =>
                           n67, ZN => n99);
   U25 : OAI22_X1 port map( A1 => net134797, A2 => n193, B1 => net134803, B2 =>
                           n60, ZN => n74);
   U26 : INV_X1 port map( A => i(28), ZN => n197);
   U27 : INV_X1 port map( A => i(27), ZN => n190);
   U28 : OAI22_X1 port map( A1 => net134801, A2 => n199, B1 => net134807, B2 =>
                           n43, ZN => n91);
   U29 : INV_X1 port map( A => i(7), ZN => n199);
   U30 : OAI22_X1 port map( A1 => net134799, A2 => n179, B1 => net134805, B2 =>
                           n50, ZN => n84);
   U31 : OAI22_X1 port map( A1 => net134799, A2 => n181, B1 => net134805, B2 =>
                           n48, ZN => n86);
   U32 : OAI22_X1 port map( A1 => n198, A2 => net134801, B1 => net134807, B2 =>
                           n36, ZN => n98);
   U33 : INV_X1 port map( A => i(0), ZN => n198);
   U34 : OAI22_X1 port map( A1 => net134799, A2 => n183, B1 => net134805, B2 =>
                           n54, ZN => n80);
   U35 : OAI22_X1 port map( A1 => n192, A2 => net134797, B1 => net134803, B2 =>
                           n61, ZN => n73);
   U36 : INV_X1 port map( A => i(17), ZN => n184);
   U37 : INV_X1 port map( A => i(12), ZN => n181);
   U38 : OAI22_X1 port map( A1 => net134797, A2 => n197, B1 => net134803, B2 =>
                           n64, ZN => n70);
   U39 : OAI22_X1 port map( A1 => net134797, A2 => n195, B1 => net134803, B2 =>
                           n66, ZN => n68);
   U40 : INV_X1 port map( A => i(16), ZN => n185);
   U41 : INV_X1 port map( A => i(13), ZN => n180);
   U42 : INV_X1 port map( A => i(5), ZN => n204);
   U43 : INV_X1 port map( A => i(24), ZN => n193);
   U44 : INV_X1 port map( A => i(14), ZN => n179);
   U45 : INV_X1 port map( A => i(9), ZN => n176);
   U46 : OAI22_X1 port map( A1 => n203, A2 => net134801, B1 => net134807, B2 =>
                           n37, ZN => n97);
   U47 : INV_X1 port map( A => i(31), ZN => n194);
   U48 : OAI22_X1 port map( A1 => net134797, A2 => n196, B1 => net134803, B2 =>
                           n65, ZN => n69);
   U49 : INV_X1 port map( A => i(15), ZN => n178);
   U50 : OAI22_X1 port map( A1 => net134799, A2 => n177, B1 => net134805, B2 =>
                           n44, ZN => n90);
   U51 : OAI22_X1 port map( A1 => net134797, A2 => n187, B1 => net134803, B2 =>
                           n58, ZN => n76);
   U52 : OAI22_X1 port map( A1 => n200, A2 => net134801, B1 => net134807, B2 =>
                           n39, ZN => n95);
   U53 : OAI22_X1 port map( A1 => net134799, A2 => n175, B1 => net134805, B2 =>
                           n46, ZN => n88);
   U54 : INV_X1 port map( A => i(18), ZN => n183);
   U55 : INV_X1 port map( A => i(21), ZN => n188);
   U56 : OAI22_X1 port map( A1 => net134797, A2 => n186, B1 => net134803, B2 =>
                           n59, ZN => n75);
   U57 : INV_X1 port map( A => i(23), ZN => n186);
   U58 : OAI22_X1 port map( A1 => n204, A2 => net134801, B1 => net134807, B2 =>
                           n41, ZN => n93);
   U59 : INV_X1 port map( A => i(3), ZN => n200);
   U60 : INV_X1 port map( A => i(30), ZN => n195);
   U61 : INV_X1 port map( A => i(26), ZN => n191);
   U62 : OAI22_X1 port map( A1 => n174, A2 => net134799, B1 => net134805, B2 =>
                           n47, ZN => n87);
   U63 : INV_X1 port map( A => i(11), ZN => n174);
   U64 : INV_X1 port map( A => i(22), ZN => n187);
   U65 : INV_X1 port map( A => i(25), ZN => n192);
   U66 : OAI22_X1 port map( A1 => n189, A2 => net134797, B1 => net134803, B2 =>
                           n56, ZN => n78);
   U67 : INV_X1 port map( A => i(20), ZN => n189);
   U68 : INV_X1 port map( A => i(8), ZN => n177);
   U69 : INV_X1 port map( A => i(6), ZN => n202);
   U70 : OAI22_X1 port map( A1 => n201, A2 => net134801, B1 => net134807, B2 =>
                           n38, ZN => n96);
   U71 : INV_X1 port map( A => i(2), ZN => n201);
   U72 : OAI22_X1 port map( A1 => net134799, A2 => n182, B1 => net134805, B2 =>
                           n55, ZN => n79);
   U73 : INV_X1 port map( A => i(19), ZN => n182);
   U74 : INV_X1 port map( A => i(1), ZN => n203);
   U75 : INV_X1 port map( A => i(29), ZN => n196);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity ALU_M32_C4 is

   port( CODE : in std_logic_vector (3 downto 0);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
         downto 0));

end ALU_M32_C4;

architecture SYN_structural of ALU_M32_C4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component COMPARATOR_M32
      port( A, B : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  OUTPUT : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4ADDER_n_bit32
      port( A, B : in std_logic_vector (31 downto 0);  cin0 : in std_logic;  S 
            : out std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_M32_N5
      port( A, B : in std_logic_vector (31 downto 0);  LEFT_RIGHT : in 
            std_logic;  OUTPUT : out std_logic_vector (31 downto 0));
   end component;
   
   signal Comparison_1_port, SHIFTERout_31_port, SHIFTERout_30_port, 
      SHIFTERout_29_port, SHIFTERout_28_port, SHIFTERout_27_port, 
      SHIFTERout_26_port, SHIFTERout_25_port, SHIFTERout_24_port, 
      SHIFTERout_23_port, SHIFTERout_22_port, SHIFTERout_21_port, 
      SHIFTERout_20_port, SHIFTERout_19_port, SHIFTERout_18_port, 
      SHIFTERout_17_port, SHIFTERout_16_port, SHIFTERout_15_port, 
      SHIFTERout_14_port, SHIFTERout_13_port, SHIFTERout_12_port, 
      SHIFTERout_11_port, SHIFTERout_10_port, SHIFTERout_9_port, 
      SHIFTERout_8_port, SHIFTERout_7_port, SHIFTERout_6_port, 
      SHIFTERout_5_port, SHIFTERout_4_port, SHIFTERout_3_port, 
      SHIFTERout_2_port, SHIFTERout_1_port, SHIFTERout_0_port, ADDERout_31_port
      , ADDERout_30_port, ADDERout_29_port, ADDERout_28_port, ADDERout_27_port,
      ADDERout_26_port, ADDERout_25_port, ADDERout_24_port, ADDERout_23_port, 
      ADDERout_22_port, ADDERout_21_port, ADDERout_20_port, ADDERout_19_port, 
      ADDERout_18_port, ADDERout_17_port, ADDERout_16_port, ADDERout_15_port, 
      ADDERout_14_port, ADDERout_13_port, ADDERout_12_port, ADDERout_11_port, 
      ADDERout_10_port, ADDERout_9_port, ADDERout_8_port, ADDERout_7_port, 
      ADDERout_6_port, ADDERout_5_port, ADDERout_4_port, ADDERout_3_port, 
      ADDERout_2_port, ADDERout_1_port, ADDERout_0_port, COMPARATORout_0_port, 
      n70, n71, n72, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n169, n170, n171, n172, net131848, net133061, 
      net134759, net134757, net134755, net134765, net134763, net134761, 
      net134777, net134775, net134773, net134771, net134769, net134767, 
      net134783, net134781, net134779, net134795, net134793, net134791, 
      net134789, net134787, net134785, net131887, net131855, n91, n90, 
      net131849, n92, n74, n73, n176, n175, n174, n173, n645, n646, n647, n648,
      n649, n650, n651, n652, n653, n654, n655, n657, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n_1030, n_1031, 
      n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, 
      n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, 
      n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, 
      n_1059, n_1060 : std_logic;

begin
   
   SHIFTOP : SHIFTER_M32_N5 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => n645, B(2) =>
                           n663, B(1) => DATA2(1), B(0) => n685, LEFT_RIGHT => 
                           CODE(0), OUTPUT(31) => SHIFTERout_31_port, 
                           OUTPUT(30) => SHIFTERout_30_port, OUTPUT(29) => 
                           SHIFTERout_29_port, OUTPUT(28) => SHIFTERout_28_port
                           , OUTPUT(27) => SHIFTERout_27_port, OUTPUT(26) => 
                           SHIFTERout_26_port, OUTPUT(25) => SHIFTERout_25_port
                           , OUTPUT(24) => SHIFTERout_24_port, OUTPUT(23) => 
                           SHIFTERout_23_port, OUTPUT(22) => SHIFTERout_22_port
                           , OUTPUT(21) => SHIFTERout_21_port, OUTPUT(20) => 
                           SHIFTERout_20_port, OUTPUT(19) => SHIFTERout_19_port
                           , OUTPUT(18) => SHIFTERout_18_port, OUTPUT(17) => 
                           SHIFTERout_17_port, OUTPUT(16) => SHIFTERout_16_port
                           , OUTPUT(15) => SHIFTERout_15_port, OUTPUT(14) => 
                           SHIFTERout_14_port, OUTPUT(13) => SHIFTERout_13_port
                           , OUTPUT(12) => SHIFTERout_12_port, OUTPUT(11) => 
                           SHIFTERout_11_port, OUTPUT(10) => SHIFTERout_10_port
                           , OUTPUT(9) => SHIFTERout_9_port, OUTPUT(8) => 
                           SHIFTERout_8_port, OUTPUT(7) => SHIFTERout_7_port, 
                           OUTPUT(6) => SHIFTERout_6_port, OUTPUT(5) => 
                           SHIFTERout_5_port, OUTPUT(4) => SHIFTERout_4_port, 
                           OUTPUT(3) => SHIFTERout_3_port, OUTPUT(2) => 
                           SHIFTERout_2_port, OUTPUT(1) => SHIFTERout_1_port, 
                           OUTPUT(0) => SHIFTERout_0_port);
   ADDSUBOP : P4ADDER_n_bit32 port map( A(31) => DATA1(31), A(30) => DATA1(30),
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => n695, B(29) => n698, B(28) => n701, B(27) 
                           => n686, B(26) => n697, B(25) => n703, B(24) => n702
                           , B(23) => n705, B(22) => n736, B(21) => n694, B(20)
                           => n688, B(19) => n691, B(18) => n708, B(17) => n711
                           , B(16) => n707, B(15) => n699, B(14) => n693, B(13)
                           => n704, B(12) => n700, B(11) => n689, B(10) => n706
                           , B(9) => n692, B(8) => n687, B(7) => n690, B(6) => 
                           n696, B(5) => DATA2(5), B(4) => DATA2(4), B(3) => 
                           DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1), B(0) 
                           => DATA2(0), cin0 => net133061, S(31) => 
                           ADDERout_31_port, S(30) => ADDERout_30_port, S(29) 
                           => ADDERout_29_port, S(28) => ADDERout_28_port, 
                           S(27) => ADDERout_27_port, S(26) => ADDERout_26_port
                           , S(25) => ADDERout_25_port, S(24) => 
                           ADDERout_24_port, S(23) => ADDERout_23_port, S(22) 
                           => ADDERout_22_port, S(21) => ADDERout_21_port, 
                           S(20) => ADDERout_20_port, S(19) => ADDERout_19_port
                           , S(18) => ADDERout_18_port, S(17) => 
                           ADDERout_17_port, S(16) => ADDERout_16_port, S(15) 
                           => ADDERout_15_port, S(14) => ADDERout_14_port, 
                           S(13) => ADDERout_13_port, S(12) => ADDERout_12_port
                           , S(11) => ADDERout_11_port, S(10) => 
                           ADDERout_10_port, S(9) => ADDERout_9_port, S(8) => 
                           ADDERout_8_port, S(7) => ADDERout_7_port, S(6) => 
                           ADDERout_6_port, S(5) => ADDERout_5_port, S(4) => 
                           ADDERout_4_port, S(3) => ADDERout_3_port, S(2) => 
                           ADDERout_2_port, S(1) => ADDERout_1_port, S(0) => 
                           ADDERout_0_port);
   COMPOP : COMPARATOR_M32 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => n695, B(29) => n698, B(28) => n701, B(27) 
                           => n686, B(26) => n697, B(25) => n703, B(24) => n702
                           , B(23) => n705, B(22) => n736, B(21) => n694, B(20)
                           => n688, B(19) => n691, B(18) => n708, B(17) => n711
                           , B(16) => n707, B(15) => n699, B(14) => n693, B(13)
                           => n704, B(12) => n700, B(11) => n689, B(10) => n706
                           , B(9) => n692, B(8) => n687, B(7) => n690, B(6) => 
                           n696, B(5) => DATA2(5), B(4) => DATA2(4), B(3) => 
                           DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1), B(0) 
                           => n685, sel(1) => Comparison_1_port, sel(0) => 
                           net131848, OUTPUT(31) => n_1030, OUTPUT(30) => 
                           n_1031, OUTPUT(29) => n_1032, OUTPUT(28) => n_1033, 
                           OUTPUT(27) => n_1034, OUTPUT(26) => n_1035, 
                           OUTPUT(25) => n_1036, OUTPUT(24) => n_1037, 
                           OUTPUT(23) => n_1038, OUTPUT(22) => n_1039, 
                           OUTPUT(21) => n_1040, OUTPUT(20) => n_1041, 
                           OUTPUT(19) => n_1042, OUTPUT(18) => n_1043, 
                           OUTPUT(17) => n_1044, OUTPUT(16) => n_1045, 
                           OUTPUT(15) => n_1046, OUTPUT(14) => n_1047, 
                           OUTPUT(13) => n_1048, OUTPUT(12) => n_1049, 
                           OUTPUT(11) => n_1050, OUTPUT(10) => n_1051, 
                           OUTPUT(9) => n_1052, OUTPUT(8) => n_1053, OUTPUT(7) 
                           => n_1054, OUTPUT(6) => n_1055, OUTPUT(5) => n_1056,
                           OUTPUT(4) => n_1057, OUTPUT(3) => n_1058, OUTPUT(2) 
                           => n_1059, OUTPUT(1) => n_1060, OUTPUT(0) => 
                           COMPARATORout_0_port);
   U209 : XOR2_X1 port map( A => CODE(1), B => CODE(0), Z => n176);
   U2 : INV_X1 port map( A => n801, ZN => n645);
   U3 : AOI221_X1 port map( B1 => net134767, B2 => n744, C1 => DATA1(30), C2 =>
                           net134781, A => net134785, ZN => n100);
   U4 : AOI221_X1 port map( B1 => net134771, B2 => n762, C1 => DATA1(12), C2 =>
                           net134779, A => net134789, ZN => n160);
   U5 : AOI221_X1 port map( B1 => net134767, B2 => n767, C1 => DATA1(7), C2 => 
                           net134783, A => net134785, ZN => n82);
   U6 : AOI221_X1 port map( B1 => net134769, B2 => n753, C1 => DATA1(21), C2 =>
                           net134781, A => net134787, ZN => n130);
   U7 : AOI221_X1 port map( B1 => net134769, B2 => n750, C1 => DATA1(24), C2 =>
                           net134781, A => net134787, ZN => n121);
   U8 : AOI221_X1 port map( B1 => net134769, B2 => n748, C1 => DATA1(26), C2 =>
                           net134781, A => net134787, ZN => n115);
   U9 : AOI221_X1 port map( B1 => net134767, B2 => n747, C1 => DATA1(27), C2 =>
                           net134781, A => net134785, ZN => n112);
   U10 : INV_X1 port map( A => CODE(0), ZN => net133061);
   U11 : NOR2_X1 port map( A1 => n90, A2 => net131887, ZN => n646);
   U12 : NOR2_X1 port map( A1 => n91, A2 => net131855, ZN => n647);
   U13 : AND2_X1 port map( A1 => n726, A2 => n725, ZN => n648);
   U14 : AND2_X1 port map( A1 => n728, A2 => n727, ZN => n649);
   U15 : AND2_X1 port map( A1 => n730, A2 => n729, ZN => n650);
   U16 : AND2_X1 port map( A1 => n714, A2 => n713, ZN => n651);
   U17 : AND2_X1 port map( A1 => n742, A2 => n741, ZN => n652);
   U18 : NOR3_X1 port map( A1 => net131848, A2 => CODE(0), A3 => n174, ZN => 
                           n77);
   U19 : NOR2_X1 port map( A1 => n130, A2 => n784, ZN => n653);
   U20 : NOR2_X1 port map( A1 => n129, A2 => n753, ZN => n654);
   U21 : NOR2_X1 port map( A1 => n653, A2 => n654, ZN => n655);
   U22 : NAND2_X1 port map( A1 => n131, A2 => n655, ZN => OUTALU(21));
   U23 : BUF_X1 port map( A => DATA2(7), Z => n690);
   U24 : BUF_X1 port map( A => DATA2(13), Z => n704);
   U25 : NOR2_X1 port map( A1 => n646, A2 => n647, ZN => n657);
   U26 : NAND2_X1 port map( A1 => n92, A2 => n657, ZN => OUTALU(4));
   U27 : OAI221_X1 port map( B1 => n659, B2 => n660, C1 => n661, C2 => n662, A 
                           => n652, ZN => OUTALU(5));
   U28 : INV_X1 port map( A => SHIFTERout_5_port, ZN => n659);
   U29 : INV_X1 port map( A => n73, ZN => n660);
   U30 : INV_X1 port map( A => ADDERout_5_port, ZN => n661);
   U31 : INV_X1 port map( A => n74, ZN => n662);
   U32 : AOI22_X1 port map( A1 => SHIFTERout_21_port, A2 => n73, B1 => 
                           ADDERout_21_port, B2 => n74, ZN => n131);
   U33 : AOI22_X1 port map( A1 => SHIFTERout_3_port, A2 => n73, B1 => 
                           ADDERout_3_port, B2 => n74, ZN => n95);
   U34 : AOI22_X1 port map( A1 => SHIFTERout_8_port, A2 => n73, B1 => 
                           ADDERout_8_port, B2 => n74, ZN => n80);
   U35 : AOI22_X1 port map( A1 => SHIFTERout_4_port, A2 => n73, B1 => 
                           ADDERout_4_port, B2 => n74, ZN => n92);
   U36 : AOI22_X1 port map( A1 => SHIFTERout_1_port, A2 => n73, B1 => 
                           ADDERout_1_port, B2 => n74, ZN => n137);
   U37 : NAND2_X1 port map( A1 => n128, A2 => n648, ZN => OUTALU(22));
   U38 : CLKBUF_X1 port map( A => DATA2(2), Z => n663);
   U39 : OR2_X1 port map( A1 => n120, A2 => n750, ZN => n664);
   U40 : OR2_X1 port map( A1 => n121, A2 => n781, ZN => n665);
   U41 : NAND3_X1 port map( A1 => n664, A2 => n665, A3 => n122, ZN => 
                           OUTALU(24));
   U42 : BUF_X1 port map( A => DATA2(15), Z => n699);
   U43 : OR2_X1 port map( A1 => n96, A2 => n743, ZN => n666);
   U44 : OR2_X1 port map( A1 => n97, A2 => n774, ZN => n667);
   U45 : NAND3_X1 port map( A1 => n98, A2 => n667, A3 => n666, ZN => OUTALU(31)
                           );
   U46 : OR2_X1 port map( A1 => n105, A2 => n745, ZN => n668);
   U47 : OR2_X1 port map( A1 => n106, A2 => n776, ZN => n669);
   U48 : NAND3_X1 port map( A1 => n107, A2 => n669, A3 => n668, ZN => 
                           OUTALU(29));
   U49 : OR2_X1 port map( A1 => n150, A2 => n759, ZN => n670);
   U50 : OR2_X1 port map( A1 => n151, A2 => n790, ZN => n671);
   U51 : NAND3_X1 port map( A1 => n670, A2 => n671, A3 => n152, ZN => 
                           OUTALU(15));
   U52 : OR2_X1 port map( A1 => n159, A2 => n762, ZN => n672);
   U53 : OR2_X1 port map( A1 => n160, A2 => n793, ZN => n673);
   U54 : NAND3_X1 port map( A1 => n161, A2 => n673, A3 => n672, ZN => 
                           OUTALU(12));
   U55 : OR2_X1 port map( A1 => n123, A2 => n751, ZN => n674);
   U56 : OR2_X1 port map( A1 => n124, A2 => n782, ZN => n675);
   U57 : NAND3_X1 port map( A1 => n674, A2 => n675, A3 => n125, ZN => 
                           OUTALU(23));
   U58 : OR2_X1 port map( A1 => n165, A2 => n764, ZN => n676);
   U59 : OR2_X1 port map( A1 => n166, A2 => n795, ZN => n677);
   U60 : NAND3_X1 port map( A1 => n676, A2 => n677, A3 => n167, ZN => 
                           OUTALU(10));
   U61 : OR2_X1 port map( A1 => n141, A2 => n756, ZN => n678);
   U62 : OR2_X1 port map( A1 => n142, A2 => n787, ZN => n679);
   U63 : NAND3_X1 port map( A1 => n143, A2 => n679, A3 => n678, ZN => 
                           OUTALU(18));
   U64 : NAND2_X1 port map( A1 => n104, A2 => n649, ZN => OUTALU(2));
   U65 : OR2_X1 port map( A1 => n78, A2 => n766, ZN => n680);
   U66 : OR2_X1 port map( A1 => n79, A2 => n797, ZN => n681);
   U67 : NAND3_X1 port map( A1 => n680, A2 => n681, A3 => n80, ZN => OUTALU(8))
                           ;
   U68 : OR2_X1 port map( A1 => n108, A2 => n746, ZN => n682);
   U69 : OR2_X1 port map( A1 => n109, A2 => n777, ZN => n683);
   U70 : NAND3_X1 port map( A1 => n682, A2 => n683, A3 => n110, ZN => 
                           OUTALU(28));
   U71 : NAND2_X1 port map( A1 => n101, A2 => n651, ZN => OUTALU(30));
   U72 : BUF_X1 port map( A => n74, Z => net134765);
   U73 : BUF_X1 port map( A => n73, Z => net134755);
   U74 : OAI21_X1 port map( B1 => Comparison_1_port, B2 => n174, A => n175, ZN 
                           => n74);
   U75 : BUF_X1 port map( A => n74, Z => net134761);
   U76 : BUF_X1 port map( A => n74, Z => net134763);
   U77 : OR3_X1 port map( A1 => CODE(2), A2 => CODE(3), A3 => n173, ZN => n175)
                           ;
   U78 : AND3_X1 port map( A1 => net131849, A2 => n684, A3 => n176, ZN => n73);
   U79 : BUF_X1 port map( A => n73, Z => net134759);
   U80 : BUF_X1 port map( A => n73, Z => net134757);
   U81 : NAND2_X1 port map( A1 => CODE(0), A2 => CODE(1), ZN => n173);
   U82 : NOR3_X1 port map( A1 => net133061, A2 => CODE(1), A3 => n174, ZN => 
                           n76);
   U83 : NAND2_X1 port map( A1 => net131848, A2 => net133061, ZN => 
                           Comparison_1_port);
   U84 : INV_X1 port map( A => CODE(3), ZN => n684);
   U85 : NAND2_X1 port map( A1 => CODE(2), A2 => n684, ZN => n174);
   U86 : INV_X1 port map( A => CODE(2), ZN => net131849);
   U87 : NAND4_X1 port map( A1 => COMPARATORout_0_port, A2 => CODE(3), A3 => 
                           n173, A4 => net131849, ZN => n172);
   U88 : NOR2_X1 port map( A1 => n174, A2 => n173, ZN => n75);
   U89 : INV_X1 port map( A => CODE(1), ZN => net131848);
   U90 : INV_X1 port map( A => DATA2(4), ZN => net131855);
   U91 : AOI21_X1 port map( B1 => net134775, B2 => net131855, A => net134793, 
                           ZN => n90);
   U92 : AOI221_X1 port map( B1 => net134767, B2 => net131887, C1 => DATA1(4), 
                           C2 => net134783, A => net134785, ZN => n91);
   U93 : BUF_X1 port map( A => n77, Z => net134785);
   U94 : BUF_X1 port map( A => n76, Z => net134783);
   U95 : INV_X1 port map( A => DATA1(4), ZN => net131887);
   U96 : BUF_X1 port map( A => n75, Z => net134767);
   U97 : BUF_X1 port map( A => n77, Z => net134793);
   U98 : BUF_X1 port map( A => n75, Z => net134775);
   U99 : INV_X1 port map( A => n804, ZN => n685);
   U100 : CLKBUF_X1 port map( A => DATA2(27), Z => n686);
   U101 : CLKBUF_X1 port map( A => DATA2(8), Z => n687);
   U102 : CLKBUF_X1 port map( A => DATA2(20), Z => n688);
   U103 : CLKBUF_X1 port map( A => DATA2(11), Z => n689);
   U104 : CLKBUF_X1 port map( A => DATA2(19), Z => n691);
   U105 : CLKBUF_X1 port map( A => DATA2(9), Z => n692);
   U106 : CLKBUF_X1 port map( A => DATA2(14), Z => n693);
   U107 : CLKBUF_X1 port map( A => DATA2(21), Z => n694);
   U108 : CLKBUF_X1 port map( A => DATA2(30), Z => n695);
   U109 : NAND2_X1 port map( A1 => n137, A2 => n650, ZN => OUTALU(1));
   U110 : CLKBUF_X1 port map( A => DATA2(6), Z => n696);
   U111 : CLKBUF_X1 port map( A => DATA2(26), Z => n697);
   U112 : CLKBUF_X1 port map( A => DATA2(29), Z => n698);
   U113 : CLKBUF_X1 port map( A => DATA2(12), Z => n700);
   U114 : CLKBUF_X1 port map( A => DATA2(28), Z => n701);
   U115 : CLKBUF_X1 port map( A => DATA2(24), Z => n702);
   U116 : CLKBUF_X1 port map( A => DATA2(25), Z => n703);
   U117 : CLKBUF_X1 port map( A => DATA2(23), Z => n705);
   U118 : CLKBUF_X1 port map( A => DATA2(10), Z => n706);
   U119 : CLKBUF_X1 port map( A => DATA2(16), Z => n707);
   U120 : CLKBUF_X1 port map( A => DATA2(18), Z => n708);
   U121 : OR2_X1 port map( A1 => n156, A2 => n761, ZN => n709);
   U122 : OR2_X1 port map( A1 => n157, A2 => n792, ZN => n710);
   U123 : NAND3_X1 port map( A1 => n158, A2 => n710, A3 => n709, ZN => 
                           OUTALU(13));
   U124 : CLKBUF_X1 port map( A => DATA2(17), Z => n711);
   U125 : NAND3_X1 port map( A1 => n733, A2 => n734, A3 => n735, ZN => 
                           OUTALU(0));
   U126 : OR2_X1 port map( A1 => n99, A2 => n744, ZN => n713);
   U127 : OR2_X1 port map( A1 => n100, A2 => n775, ZN => n714);
   U128 : OR2_X1 port map( A1 => n70, A2 => n765, ZN => n715);
   U129 : OR2_X1 port map( A1 => n71, A2 => n796, ZN => n716);
   U130 : NAND3_X1 port map( A1 => n72, A2 => n716, A3 => n715, ZN => OUTALU(9)
                           );
   U131 : OR2_X1 port map( A1 => n144, A2 => n757, ZN => n717);
   U132 : OR2_X1 port map( A1 => n145, A2 => n788, ZN => n718);
   U133 : NAND3_X1 port map( A1 => n717, A2 => n718, A3 => n146, ZN => 
                           OUTALU(17));
   U134 : OR2_X1 port map( A1 => n93, A2 => n770, ZN => n719);
   U135 : OR2_X1 port map( A1 => n94, A2 => n801, ZN => n720);
   U136 : NAND3_X1 port map( A1 => n95, A2 => n720, A3 => n719, ZN => OUTALU(3)
                           );
   U137 : OR2_X1 port map( A1 => n117, A2 => n749, ZN => n721);
   U138 : OR2_X1 port map( A1 => n118, A2 => n780, ZN => n722);
   U139 : NAND3_X1 port map( A1 => n119, A2 => n722, A3 => n721, ZN => 
                           OUTALU(25));
   U140 : OR2_X1 port map( A1 => n162, A2 => n763, ZN => n723);
   U141 : OR2_X1 port map( A1 => n163, A2 => n794, ZN => n724);
   U142 : NAND3_X1 port map( A1 => n164, A2 => n724, A3 => n723, ZN => 
                           OUTALU(11));
   U143 : OR2_X1 port map( A1 => n126, A2 => n752, ZN => n725);
   U144 : OR2_X1 port map( A1 => n127, A2 => n783, ZN => n726);
   U145 : OR2_X1 port map( A1 => n102, A2 => n771, ZN => n727);
   U146 : OR2_X1 port map( A1 => n103, A2 => n802, ZN => n728);
   U147 : OR2_X1 port map( A1 => n135, A2 => n772, ZN => n729);
   U148 : OR2_X1 port map( A1 => n136, A2 => n803, ZN => n730);
   U149 : OR2_X1 port map( A1 => n84, A2 => n768, ZN => n731);
   U150 : OR2_X1 port map( A1 => n85, A2 => n799, ZN => n732);
   U151 : NAND3_X1 port map( A1 => n86, A2 => n732, A3 => n731, ZN => OUTALU(6)
                           );
   U152 : NAND2_X1 port map( A1 => SHIFTERout_0_port, A2 => net134759, ZN => 
                           n733);
   U153 : NAND2_X1 port map( A1 => ADDERout_0_port, A2 => net134761, ZN => n734
                           );
   U154 : INV_X1 port map( A => n169, ZN => n735);
   U155 : BUF_X1 port map( A => n75, Z => net134771);
   U156 : BUF_X1 port map( A => n75, Z => net134769);
   U157 : BUF_X1 port map( A => n75, Z => net134773);
   U158 : BUF_X1 port map( A => n77, Z => net134789);
   U159 : BUF_X1 port map( A => n77, Z => net134791);
   U160 : BUF_X1 port map( A => n77, Z => net134787);
   U161 : AOI22_X1 port map( A1 => SHIFTERout_14_port, A2 => net134759, B1 => 
                           ADDERout_14_port, B2 => net134761, ZN => n155);
   U162 : AOI22_X1 port map( A1 => SHIFTERout_15_port, A2 => net134759, B1 => 
                           ADDERout_15_port, B2 => net134761, ZN => n152);
   U163 : AOI22_X1 port map( A1 => SHIFTERout_10_port, A2 => net134759, B1 => 
                           ADDERout_10_port, B2 => net134761, ZN => n167);
   U164 : AOI22_X1 port map( A1 => SHIFTERout_19_port, A2 => net134757, B1 => 
                           ADDERout_19_port, B2 => net134761, ZN => n140);
   U165 : AOI221_X1 port map( B1 => net134769, B2 => n755, C1 => DATA1(19), C2 
                           => net134779, A => net134787, ZN => n139);
   U166 : AOI221_X1 port map( B1 => net134767, B2 => n746, C1 => DATA1(28), C2 
                           => net134781, A => net134785, ZN => n109);
   U167 : AOI221_X1 port map( B1 => net134769, B2 => n765, C1 => net134783, C2 
                           => DATA1(9), A => net134787, ZN => n71);
   U168 : AOI221_X1 port map( B1 => net134769, B2 => n772, C1 => DATA1(1), C2 
                           => net134779, A => net134787, ZN => n136);
   U169 : AOI221_X1 port map( B1 => net134771, B2 => n761, C1 => DATA1(13), C2 
                           => net134779, A => net134789, ZN => n157);
   U170 : AOI221_X1 port map( B1 => net134767, B2 => n770, C1 => DATA1(3), C2 
                           => net134783, A => net134785, ZN => n94);
   U171 : AOI221_X1 port map( B1 => net134769, B2 => n749, C1 => DATA1(25), C2 
                           => net134781, A => net134787, ZN => n118);
   U172 : AOI221_X1 port map( B1 => net134769, B2 => n751, C1 => DATA1(23), C2 
                           => net134781, A => net134787, ZN => n124);
   U173 : AOI221_X1 port map( B1 => net134767, B2 => n768, C1 => DATA1(6), C2 
                           => net134783, A => net134785, ZN => n85);
   U174 : AOI221_X1 port map( B1 => net134767, B2 => n766, C1 => DATA1(8), C2 
                           => net134783, A => net134785, ZN => n79);
   U175 : AOI221_X1 port map( B1 => net134771, B2 => n763, C1 => DATA1(11), C2 
                           => net134779, A => net134789, ZN => n163);
   U176 : AOI221_X1 port map( B1 => net134771, B2 => n760, C1 => DATA1(14), C2 
                           => net134779, A => net134789, ZN => n154);
   U177 : AOI221_X1 port map( B1 => net134771, B2 => n759, C1 => DATA1(15), C2 
                           => net134779, A => net134789, ZN => n151);
   U178 : AOI221_X1 port map( B1 => net134771, B2 => n757, C1 => DATA1(17), C2 
                           => net134779, A => net134789, ZN => n145);
   U179 : AOI221_X1 port map( B1 => net134769, B2 => n756, C1 => DATA1(18), C2 
                           => net134779, A => net134787, ZN => n142);
   U180 : AOI221_X1 port map( B1 => net134769, B2 => n752, C1 => DATA1(22), C2 
                           => net134781, A => net134787, ZN => n127);
   U181 : AOI221_X1 port map( B1 => net134767, B2 => n745, C1 => DATA1(29), C2 
                           => net134781, A => net134785, ZN => n106);
   U182 : AOI221_X1 port map( B1 => net134767, B2 => n743, C1 => DATA1(31), C2 
                           => net134783, A => net134785, ZN => n97);
   U183 : BUF_X1 port map( A => n76, Z => net134779);
   U184 : BUF_X1 port map( A => n76, Z => net134781);
   U185 : INV_X1 port map( A => DATA1(30), ZN => n744);
   U186 : INV_X1 port map( A => DATA1(29), ZN => n745);
   U187 : INV_X1 port map( A => DATA1(25), ZN => n749);
   U188 : INV_X1 port map( A => DATA1(1), ZN => n772);
   U189 : INV_X1 port map( A => DATA1(22), ZN => n752);
   U190 : INV_X1 port map( A => DATA1(26), ZN => n748);
   U191 : INV_X1 port map( A => DATA1(23), ZN => n751);
   U192 : INV_X1 port map( A => DATA1(31), ZN => n743);
   U193 : INV_X1 port map( A => DATA1(28), ZN => n746);
   U194 : INV_X1 port map( A => DATA1(13), ZN => n761);
   U195 : INV_X1 port map( A => DATA1(8), ZN => n766);
   U196 : INV_X1 port map( A => DATA1(19), ZN => n755);
   U197 : INV_X1 port map( A => DATA1(6), ZN => n768);
   U198 : INV_X1 port map( A => DATA1(15), ZN => n759);
   U199 : INV_X1 port map( A => DATA1(17), ZN => n757);
   U200 : INV_X1 port map( A => DATA1(18), ZN => n756);
   U201 : INV_X1 port map( A => DATA1(21), ZN => n753);
   U202 : INV_X1 port map( A => DATA1(24), ZN => n750);
   U203 : INV_X1 port map( A => DATA1(12), ZN => n762);
   U204 : INV_X1 port map( A => DATA1(7), ZN => n767);
   U205 : INV_X1 port map( A => DATA1(14), ZN => n760);
   U206 : INV_X1 port map( A => DATA1(27), ZN => n747);
   U207 : INV_X1 port map( A => DATA1(9), ZN => n765);
   U208 : INV_X1 port map( A => DATA1(11), ZN => n763);
   U210 : INV_X1 port map( A => DATA1(3), ZN => n770);
   U211 : INV_X1 port map( A => DATA1(0), ZN => n773);
   U212 : INV_X1 port map( A => n711, ZN => n788);
   U213 : INV_X1 port map( A => n687, ZN => n797);
   U214 : INV_X1 port map( A => n686, ZN => n778);
   U215 : INV_X1 port map( A => n697, ZN => n779);
   U216 : INV_X1 port map( A => DATA2(1), ZN => n803);
   U217 : INV_X1 port map( A => n663, ZN => n802);
   U218 : INV_X1 port map( A => DATA2(3), ZN => n801);
   U219 : AOI221_X1 port map( B1 => net134769, B2 => n758, C1 => DATA1(16), C2 
                           => net134779, A => net134787, ZN => n148);
   U220 : AOI221_X1 port map( B1 => net134769, B2 => n754, C1 => DATA1(20), C2 
                           => net134781, A => net134787, ZN => n133);
   U221 : AOI221_X1 port map( B1 => net134767, B2 => n769, C1 => DATA1(5), C2 
                           => net134783, A => net134785, ZN => n88);
   U222 : AOI221_X1 port map( B1 => net134767, B2 => n771, C1 => DATA1(2), C2 
                           => net134781, A => net134785, ZN => n103);
   U223 : AOI221_X1 port map( B1 => net134771, B2 => n764, C1 => DATA1(10), C2 
                           => net134779, A => net134789, ZN => n166);
   U224 : AOI21_X1 port map( B1 => net134777, B2 => n804, A => net134795, ZN =>
                           n170);
   U225 : AOI221_X1 port map( B1 => net134771, B2 => n773, C1 => DATA1(0), C2 
                           => net134779, A => net134789, ZN => n171);
   U226 : AOI21_X1 port map( B1 => net134773, B2 => n778, A => net134791, ZN =>
                           n111);
   U227 : AOI21_X1 port map( B1 => net134773, B2 => n791, A => net134791, ZN =>
                           n153);
   U228 : AOI21_X1 port map( B1 => net134771, B2 => n783, A => net134789, ZN =>
                           n126);
   U229 : AOI21_X1 port map( B1 => net134771, B2 => n786, A => net134789, ZN =>
                           n138);
   U230 : AOI21_X1 port map( B1 => net134773, B2 => n782, A => net134791, ZN =>
                           n123);
   U231 : AOI21_X1 port map( B1 => net134773, B2 => n787, A => net134791, ZN =>
                           n141);
   U232 : AOI21_X1 port map( B1 => net134773, B2 => n780, A => net134791, ZN =>
                           n117);
   U233 : AOI21_X1 port map( B1 => net134773, B2 => n777, A => net134791, ZN =>
                           n108);
   U234 : AOI21_X1 port map( B1 => net134775, B2 => n792, A => net134793, ZN =>
                           n156);
   U235 : AOI21_X1 port map( B1 => net134773, B2 => n788, A => net134791, ZN =>
                           n144);
   U236 : AOI21_X1 port map( B1 => net134773, B2 => n779, A => net134791, ZN =>
                           n114);
   U237 : AOI21_X1 port map( B1 => net134775, B2 => n776, A => net134793, ZN =>
                           n105);
   U238 : AOI21_X1 port map( B1 => net134775, B2 => n775, A => net134793, ZN =>
                           n99);
   U239 : AOI21_X1 port map( B1 => net134771, B2 => n784, A => net134789, ZN =>
                           n129);
   U240 : AOI21_X1 port map( B1 => net134775, B2 => n794, A => net134793, ZN =>
                           n162);
   U241 : AOI21_X1 port map( B1 => net134777, B2 => n796, A => net134795, ZN =>
                           n70);
   U242 : AOI21_X1 port map( B1 => net134775, B2 => n799, A => net134793, ZN =>
                           n84);
   U243 : AOI21_X1 port map( B1 => net134773, B2 => n781, A => net134791, ZN =>
                           n120);
   U244 : AOI21_X1 port map( B1 => net134777, B2 => n797, A => net134793, ZN =>
                           n78);
   U245 : AOI21_X1 port map( B1 => net134775, B2 => n793, A => net134793, ZN =>
                           n159);
   U246 : AOI21_X1 port map( B1 => net134775, B2 => n801, A => net134793, ZN =>
                           n93);
   U247 : AOI21_X1 port map( B1 => net134775, B2 => n798, A => net134793, ZN =>
                           n81);
   U248 : AOI21_X1 port map( B1 => net134775, B2 => n774, A => net134793, ZN =>
                           n96);
   U249 : AOI21_X1 port map( B1 => net134773, B2 => n802, A => net134791, ZN =>
                           n102);
   U250 : AOI21_X1 port map( B1 => net134771, B2 => n803, A => net134789, ZN =>
                           n135);
   U251 : AOI21_X1 port map( B1 => net134775, B2 => n790, A => net134791, ZN =>
                           n150);
   U252 : AOI21_X1 port map( B1 => net134777, B2 => n795, A => net134793, ZN =>
                           n165);
   U253 : INV_X1 port map( A => DATA1(2), ZN => n771);
   U254 : INV_X1 port map( A => DATA1(10), ZN => n764);
   U255 : INV_X1 port map( A => n693, ZN => n791);
   U256 : INV_X1 port map( A => n704, ZN => n792);
   U257 : INV_X1 port map( A => n700, ZN => n793);
   U258 : AOI22_X1 port map( A1 => SHIFTERout_26_port, A2 => net134757, B1 => 
                           ADDERout_26_port, B2 => net134763, ZN => n116);
   U259 : INV_X1 port map( A => n695, ZN => n775);
   U260 : AOI22_X1 port map( A1 => SHIFTERout_18_port, A2 => net134757, B1 => 
                           ADDERout_18_port, B2 => net134761, ZN => n143);
   U261 : OAI221_X1 port map( B1 => n170, B2 => n773, C1 => n171, C2 => n804, A
                           => n172, ZN => n169);
   U262 : AOI22_X1 port map( A1 => SHIFTERout_24_port, A2 => net134757, B1 => 
                           ADDERout_24_port, B2 => net134763, ZN => n122);
   U263 : AOI22_X1 port map( A1 => SHIFTERout_31_port, A2 => net134755, B1 => 
                           ADDERout_31_port, B2 => net134765, ZN => n98);
   U264 : CLKBUF_X1 port map( A => DATA2(22), Z => n736);
   U265 : OR2_X1 port map( A1 => n147, A2 => n758, ZN => n737);
   U266 : OR2_X1 port map( A1 => n148, A2 => n789, ZN => n738);
   U267 : NAND3_X1 port map( A1 => n149, A2 => n738, A3 => n737, ZN => 
                           OUTALU(16));
   U268 : AOI21_X1 port map( B1 => net134773, B2 => n789, A => net134791, ZN =>
                           n147);
   U269 : INV_X1 port map( A => DATA1(16), ZN => n758);
   U270 : AOI22_X1 port map( A1 => SHIFTERout_11_port, A2 => net134759, B1 => 
                           ADDERout_11_port, B2 => net134761, ZN => n164);
   U271 : OR2_X1 port map( A1 => n132, A2 => n754, ZN => n739);
   U272 : OR2_X1 port map( A1 => n133, A2 => n785, ZN => n740);
   U273 : NAND3_X1 port map( A1 => n739, A2 => n740, A3 => n134, ZN => 
                           OUTALU(20));
   U274 : AOI21_X1 port map( B1 => net134773, B2 => n785, A => net134791, ZN =>
                           n132);
   U275 : INV_X1 port map( A => DATA1(20), ZN => n754);
   U276 : AOI22_X1 port map( A1 => SHIFTERout_25_port, A2 => net134757, B1 => 
                           ADDERout_25_port, B2 => net134763, ZN => n119);
   U277 : AOI22_X1 port map( A1 => SHIFTERout_22_port, A2 => net134757, B1 => 
                           ADDERout_22_port, B2 => net134763, ZN => n128);
   U278 : AOI22_X1 port map( A1 => SHIFTERout_23_port, A2 => net134757, B1 => 
                           ADDERout_23_port, B2 => net134763, ZN => n125);
   U279 : AOI22_X1 port map( A1 => SHIFTERout_9_port, A2 => net134755, B1 => 
                           ADDERout_9_port, B2 => net134765, ZN => n72);
   U280 : INV_X1 port map( A => n698, ZN => n776);
   U281 : INV_X1 port map( A => n708, ZN => n787);
   U282 : OAI221_X1 port map( B1 => n138, B2 => n755, C1 => n139, C2 => n786, A
                           => n140, ZN => OUTALU(19));
   U283 : AOI22_X1 port map( A1 => SHIFTERout_17_port, A2 => net134757, B1 => 
                           ADDERout_17_port, B2 => net134761, ZN => n146);
   U284 : OR2_X1 port map( A1 => n87, A2 => n769, ZN => n741);
   U285 : OR2_X1 port map( A1 => n88, A2 => n800, ZN => n742);
   U286 : AOI21_X1 port map( B1 => net134775, B2 => n800, A => net134793, ZN =>
                           n87);
   U287 : INV_X1 port map( A => DATA1(5), ZN => n769);
   U288 : INV_X1 port map( A => DATA2(5), ZN => n800);
   U289 : INV_X1 port map( A => n692, ZN => n796);
   U290 : AOI22_X1 port map( A1 => SHIFTERout_16_port, A2 => net134759, B1 => 
                           ADDERout_16_port, B2 => net134761, ZN => n149);
   U291 : INV_X1 port map( A => n691, ZN => n786);
   U292 : AOI22_X1 port map( A1 => SHIFTERout_20_port, A2 => net134757, B1 => 
                           ADDERout_20_port, B2 => net134763, ZN => n134);
   U293 : INV_X1 port map( A => DATA2(31), ZN => n774);
   U294 : OAI221_X1 port map( B1 => n153, B2 => n760, C1 => n154, C2 => n791, A
                           => n155, ZN => OUTALU(14));
   U295 : INV_X1 port map( A => n690, ZN => n798);
   U296 : AOI22_X1 port map( A1 => SHIFTERout_6_port, A2 => net134755, B1 => 
                           ADDERout_6_port, B2 => net134765, ZN => n86);
   U297 : AOI22_X1 port map( A1 => SHIFTERout_30_port, A2 => net134755, B1 => 
                           ADDERout_30_port, B2 => net134763, ZN => n101);
   U298 : INV_X1 port map( A => n694, ZN => n784);
   U299 : AOI22_X1 port map( A1 => SHIFTERout_13_port, A2 => net134759, B1 => 
                           ADDERout_13_port, B2 => net134761, ZN => n158);
   U300 : AOI22_X1 port map( A1 => SHIFTERout_12_port, A2 => net134759, B1 => 
                           ADDERout_12_port, B2 => net134761, ZN => n161);
   U301 : AOI22_X1 port map( A1 => SHIFTERout_2_port, A2 => net134755, B1 => 
                           ADDERout_2_port, B2 => net134763, ZN => n104);
   U302 : INV_X1 port map( A => n699, ZN => n790);
   U303 : OAI221_X1 port map( B1 => n81, B2 => n767, C1 => n82, C2 => n798, A 
                           => n83, ZN => OUTALU(7));
   U304 : AOI22_X1 port map( A1 => SHIFTERout_7_port, A2 => net134755, B1 => 
                           ADDERout_7_port, B2 => net134765, ZN => n83);
   U305 : INV_X1 port map( A => DATA2(0), ZN => n804);
   U306 : AOI22_X1 port map( A1 => SHIFTERout_29_port, A2 => net134755, B1 => 
                           ADDERout_29_port, B2 => net134763, ZN => n107);
   U307 : INV_X1 port map( A => n707, ZN => n789);
   U308 : INV_X1 port map( A => n688, ZN => n785);
   U309 : INV_X1 port map( A => n703, ZN => n780);
   U310 : OAI221_X1 port map( B1 => n114, B2 => n748, C1 => n115, C2 => n779, A
                           => n116, ZN => OUTALU(26));
   U311 : INV_X1 port map( A => n689, ZN => n794);
   U312 : INV_X1 port map( A => n705, ZN => n782);
   U313 : INV_X1 port map( A => n702, ZN => n781);
   U314 : AOI22_X1 port map( A1 => SHIFTERout_27_port, A2 => net134757, B1 => 
                           ADDERout_27_port, B2 => net134763, ZN => n113);
   U315 : OAI221_X1 port map( B1 => n111, B2 => n747, C1 => n112, C2 => n778, A
                           => n113, ZN => OUTALU(27));
   U316 : INV_X1 port map( A => n706, ZN => n795);
   U317 : INV_X1 port map( A => n696, ZN => n799);
   U318 : INV_X1 port map( A => n701, ZN => n777);
   U319 : AOI22_X1 port map( A1 => SHIFTERout_28_port, A2 => net134755, B1 => 
                           ADDERout_28_port, B2 => net134763, ZN => n110);
   U320 : INV_X1 port map( A => n736, ZN => n783);
   U321 : CLKBUF_X1 port map( A => n77, Z => net134795);
   U322 : CLKBUF_X1 port map( A => n75, Z => net134777);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Mux21_4 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end Mux21_4;

architecture SYN_Behavioral of Mux21_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, net133025, net133017, net133015, net133013, net133009, net133005, 
      net133003, net133001, net141441, net141472, net141479, net141488, 
      net141492, net141590, n42, n172, n173, n174, n175, n177, n178 : std_logic
      ;

begin
   
   U1 : CLKBUF_X1 port map( A => net133009, Z => net141590);
   U2 : CLKBUF_X1 port map( A => net141441, Z => n172);
   U3 : AOI22_X1 port map( A1 => net141479, A2 => a(30), B1 => net133009, B2 =>
                           b(30), ZN => n42);
   U4 : INV_X1 port map( A => n42, ZN => y(30));
   U5 : BUF_X1 port map( A => n174, Z => n173);
   U6 : AOI22_X1 port map( A1 => net133003, A2 => a(12), B1 => n173, B2 => 
                           b(12), ZN => n62);
   U7 : AOI22_X1 port map( A1 => net141492, A2 => a(11), B1 => n173, B2 => 
                           b(11), ZN => n63);
   U8 : AOI22_X1 port map( A1 => net133001, A2 => a(10), B1 => net133017, B2 =>
                           b(10), ZN => n64);
   U9 : INV_X1 port map( A => sel, ZN => n174);
   U10 : BUF_X1 port map( A => n174, Z => net133005);
   U11 : INV_X1 port map( A => n174, ZN => net133003);
   U12 : INV_X1 port map( A => n174, ZN => net141492);
   U13 : INV_X1 port map( A => n175, ZN => net141479);
   U14 : INV_X1 port map( A => sel, ZN => n175);
   U15 : BUF_X2 port map( A => n175, Z => net133009);
   U16 : BUF_X2 port map( A => n175, Z => net133017);
   U17 : INV_X1 port map( A => sel, ZN => net133025);
   U18 : CLKBUF_X1 port map( A => net141441, Z => net141488);
   U19 : BUF_X1 port map( A => net133025, Z => net133015);
   U20 : INV_X1 port map( A => net133025, ZN => net133001);
   U21 : INV_X1 port map( A => net133003, ZN => net141472);
   U22 : INV_X1 port map( A => net133025, ZN => net141441);
   U23 : OR2_X1 port map( A1 => n177, A2 => n178, ZN => y(28));
   U24 : AND2_X1 port map( A1 => net133001, A2 => a(28), ZN => n177);
   U25 : AND2_X1 port map( A1 => net133009, A2 => b(28), ZN => n178);
   U26 : BUF_X1 port map( A => net133025, Z => net133013);
   U27 : INV_X1 port map( A => n43, ZN => y(2));
   U28 : INV_X1 port map( A => n54, ZN => y(1));
   U29 : INV_X1 port map( A => n40, ZN => y(3));
   U30 : INV_X1 port map( A => n39, ZN => y(4));
   U31 : INV_X1 port map( A => n38, ZN => y(5));
   U32 : AOI22_X1 port map( A1 => a(4), A2 => net141488, B1 => b(4), B2 => 
                           net141472, ZN => n39);
   U33 : AOI22_X1 port map( A1 => a(5), A2 => net141441, B1 => b(5), B2 => 
                           net141590, ZN => n38);
   U34 : AOI22_X1 port map( A1 => a(3), A2 => n172, B1 => b(3), B2 => net141472
                           , ZN => n40);
   U35 : AOI22_X1 port map( A1 => net141479, A2 => a(9), B1 => n173, B2 => b(9)
                           , ZN => n34);
   U36 : INV_X1 port map( A => n36, ZN => y(7));
   U37 : AOI22_X1 port map( A1 => a(7), A2 => net133003, B1 => b(7), B2 => 
                           net133013, ZN => n36);
   U38 : INV_X1 port map( A => n34, ZN => y(9));
   U39 : AOI22_X1 port map( A1 => a(6), A2 => net141441, B1 => net133005, B2 =>
                           b(6), ZN => n37);
   U40 : INV_X1 port map( A => n57, ZN => y(17));
   U41 : INV_X1 port map( A => n46, ZN => y(27));
   U42 : INV_X1 port map( A => n52, ZN => y(21));
   U43 : INV_X1 port map( A => n56, ZN => y(18));
   U44 : INV_X1 port map( A => n47, ZN => y(26));
   U45 : INV_X1 port map( A => n55, ZN => y(19));
   U46 : INV_X1 port map( A => n59, ZN => y(15));
   U47 : INV_X1 port map( A => n44, ZN => y(29));
   U48 : INV_X1 port map( A => n65, ZN => y(0));
   U49 : INV_X1 port map( A => n35, ZN => y(8));
   U50 : AOI22_X1 port map( A1 => a(8), A2 => net133003, B1 => b(8), B2 => 
                           net133005, ZN => n35);
   U51 : INV_X1 port map( A => n58, ZN => y(16));
   U52 : INV_X1 port map( A => n53, ZN => y(20));
   U53 : INV_X1 port map( A => n63, ZN => y(11));
   U54 : INV_X1 port map( A => n37, ZN => y(6));
   U55 : INV_X1 port map( A => n60, ZN => y(14));
   U56 : INV_X1 port map( A => n41, ZN => y(31));
   U57 : INV_X1 port map( A => n48, ZN => y(25));
   U58 : INV_X1 port map( A => n62, ZN => y(12));
   U59 : INV_X1 port map( A => n49, ZN => y(24));
   U60 : INV_X1 port map( A => n50, ZN => y(23));
   U61 : AOI22_X1 port map( A1 => a(31), A2 => net141441, B1 => net133005, B2 
                           => b(31), ZN => n41);
   U62 : INV_X1 port map( A => n61, ZN => y(13));
   U63 : AOI22_X1 port map( A1 => a(2), A2 => net141488, B1 => b(2), B2 => 
                           net141472, ZN => n43);
   U64 : INV_X1 port map( A => n51, ZN => y(22));
   U65 : AOI22_X1 port map( A1 => net133003, A2 => a(27), B1 => net133013, B2 
                           => b(27), ZN => n46);
   U66 : AOI22_X1 port map( A1 => a(26), A2 => net141479, B1 => b(26), B2 => 
                           net133017, ZN => n47);
   U67 : AOI22_X1 port map( A1 => net133001, A2 => a(29), B1 => net133015, B2 
                           => b(29), ZN => n44);
   U68 : AOI22_X1 port map( A1 => a(20), A2 => net133003, B1 => b(20), B2 => 
                           net133017, ZN => n53);
   U69 : AOI22_X1 port map( A1 => net141479, A2 => a(21), B1 => net133013, B2 
                           => b(21), ZN => n52);
   U70 : AOI22_X1 port map( A1 => net141479, A2 => a(25), B1 => net133009, B2 
                           => b(25), ZN => n48);
   U71 : AOI22_X1 port map( A1 => net133001, A2 => a(24), B1 => net133009, B2 
                           => b(24), ZN => n49);
   U72 : AOI22_X1 port map( A1 => net141479, A2 => a(23), B1 => net133009, B2 
                           => b(23), ZN => n50);
   U73 : AOI22_X1 port map( A1 => net133001, A2 => a(22), B1 => net133015, B2 
                           => b(22), ZN => n51);
   U74 : AOI22_X1 port map( A1 => a(1), A2 => net141441, B1 => net141590, B2 =>
                           b(1), ZN => n54);
   U75 : AOI22_X1 port map( A1 => a(0), A2 => net141441, B1 => b(0), B2 => 
                           net133017, ZN => n65);
   U76 : INV_X1 port map( A => n64, ZN => y(10));
   U77 : AOI22_X1 port map( A1 => net141492, A2 => a(19), B1 => n173, B2 => 
                           b(19), ZN => n55);
   U78 : AOI22_X1 port map( A1 => net141492, A2 => a(18), B1 => net133015, B2 
                           => b(18), ZN => n56);
   U79 : AOI22_X1 port map( A1 => a(17), A2 => net141492, B1 => net133013, B2 
                           => b(17), ZN => n57);
   U80 : AOI22_X1 port map( A1 => a(14), A2 => net133003, B1 => b(14), B2 => 
                           net133017, ZN => n60);
   U81 : AOI22_X1 port map( A1 => net141492, A2 => a(16), B1 => net133005, B2 
                           => b(16), ZN => n58);
   U82 : AOI22_X1 port map( A1 => net141441, A2 => a(15), B1 => net133005, B2 
                           => b(15), ZN => n59);
   U83 : AOI22_X1 port map( A1 => net141492, A2 => a(13), B1 => b(13), B2 => 
                           net133017, ZN => n61);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity DecodeUnit_DW01_add_0 is

   port( A, B : in std_logic_vector (9 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (9 downto 0);  CO : out std_logic);

end DecodeUnit_DW01_add_0;

architecture SYN_rpl of DecodeUnit_DW01_add_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port,
      carry_4_port, carry_3_port, carry_2_port, n2, n3, n4, n5, n6, n7, n8, n9,
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19 : std_logic;

begin
   
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U3 : XOR2_X1 port map( A => A(6), B => B(6), Z => n3);
   U4 : XOR2_X1 port map( A => n3, B => carry_6_port, Z => SUM(6));
   U8 : NAND3_X1 port map( A1 => n4, A2 => n5, A3 => n6, ZN => carry_7_port);
   U9 : XOR2_X1 port map( A => A(7), B => B(7), Z => n7);
   U10 : XOR2_X1 port map( A => n7, B => carry_7_port, Z => SUM(7));
   U14 : NAND3_X1 port map( A1 => n8, A2 => n9, A3 => n10, ZN => carry_8_port);
   U15 : XOR2_X1 port map( A => B(1), B => A(1), Z => n11);
   U16 : XOR2_X1 port map( A => n2, B => n11, Z => SUM(1));
   U20 : NAND3_X1 port map( A1 => n12, A2 => n13, A3 => n14, ZN => carry_2_port
                           );
   U21 : XOR2_X1 port map( A => B(2), B => A(2), Z => n15);
   U22 : XOR2_X1 port map( A => carry_2_port, B => n15, Z => SUM(2));
   U26 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => n18, ZN => carry_3_port
                           );
   U27 : XOR2_X1 port map( A => B(9), B => A(9), Z => n19);
   U28 : XOR2_X1 port map( A => carry_9_port, B => n19, Z => SUM(9));
   U2 : NAND2_X1 port map( A1 => B(7), A2 => carry_7_port, ZN => n10);
   U5 : NAND2_X1 port map( A1 => A(6), A2 => B(6), ZN => n4);
   U6 : NAND2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => n5);
   U7 : NAND2_X1 port map( A1 => B(6), A2 => carry_6_port, ZN => n6);
   U11 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n14);
   U12 : NAND2_X1 port map( A1 => n2, A2 => B(1), ZN => n12);
   U13 : NAND2_X1 port map( A1 => n2, A2 => A(1), ZN => n13);
   U17 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => n18);
   U18 : NAND2_X1 port map( A1 => carry_2_port, A2 => B(2), ZN => n16);
   U19 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);
   U23 : NAND2_X1 port map( A1 => A(7), A2 => B(7), ZN => n8);
   U24 : NAND2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => n9);
   U25 : NAND2_X1 port map( A1 => carry_2_port, A2 => A(2), ZN => n17);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity register_file is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file;

architecture SYN_A of register_file is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
      n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, 
      n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, 
      n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, 
      n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
      n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
      n3002, n3003, n3004, n3005, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
      n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
      n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
      n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
      n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
      n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
      n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, 
      n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
      n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, 
      n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
      n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, 
      n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, 
      n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, 
      n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, 
      n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
      n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
      n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
      n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, 
      n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, 
      n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, 
      n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, 
      n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, 
      n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, 
      n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, 
      n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, 
      n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, 
      n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, 
      n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3448, n3450, 
      n3452, n3453, n3456, n3458, n3459, n3460, n3461, n3462, n3464, n3466, 
      n3468, n3469, n3472, n3474, n3475, n3476, n3477, n3478, n3480, n3482, 
      n3484, n3485, n3488, n3490, n3491, n3492, n3493, n3494, n3496, n3498, 
      n3500, n3501, n3504, n3506, n3507, n3508, n3509, n3510, n3512, n3514, 
      n3516, n3517, n3520, n3522, n3523, n3524, n3525, n3526, n3528, n3530, 
      n3532, n3533, n3536, n3538, n3539, n3540, n3541, n3542, n3544, n3546, 
      n3548, n3549, n3552, n3554, n3555, n3556, n3557, n3558, n3560, n3562, 
      n3564, n3565, n3568, n3570, n3571, n3572, n3573, n3574, n3576, n3578, 
      n3580, n3581, n3584, n3586, n3587, n3588, n3589, n3590, n3592, n3594, 
      n3596, n3597, n3600, n3602, n3603, n3604, n3605, n3606, n3608, n3610, 
      n3612, n3613, n3616, n3618, n3619, n3620, n3621, n3622, n3624, n3626, 
      n3628, n3629, n3632, n3634, n3635, n3636, n3637, n3638, n3640, n3642, 
      n3644, n3645, n3648, n3650, n3651, n3652, n3653, n3654, n3656, n3658, 
      n3660, n3661, n3664, n3666, n3667, n3668, n3669, n3670, n3672, n3674, 
      n3676, n3677, n3680, n3682, n3683, n3684, n3685, n3686, n3688, n3690, 
      n3692, n3693, n3696, n3698, n3699, n3700, n3701, n3702, n3704, n3706, 
      n3708, n3709, n3712, n3714, n3715, n3716, n3717, n3718, n3720, n3722, 
      n3724, n3725, n3728, n3730, n3731, n3732, n3733, n3734, n3736, n3738, 
      n3740, n3741, n3744, n3746, n3747, n3748, n3749, n3750, n3752, n3754, 
      n3756, n3757, n3760, n3762, n3763, n3764, n3765, n3766, n3768, n3770, 
      n3772, n3773, n3776, n3778, n3779, n3780, n3781, n3782, n3784, n3786, 
      n3788, n3789, n3792, n3794, n3795, n3796, n3797, n3798, n3800, n3802, 
      n3804, n3805, n3808, n3810, n3811, n3812, n3813, n3814, n3816, n3818, 
      n3820, n3821, n3824, n3826, n3827, n3828, n3829, n3830, n3832, n3834, 
      n3836, n3837, n3840, n3842, n3843, n3844, n3845, n3846, n3848, n3850, 
      n3852, n3853, n3856, n3858, n3859, n3860, n3861, n3862, n3864, n3866, 
      n3868, n3869, n3872, n3874, n3875, n3876, n3877, n3878, n3880, n3882, 
      n3884, n3885, n3888, n3890, n3891, n3892, n3893, n3894, n3896, n3898, 
      n3900, n3901, n3904, n3906, n3907, n3908, n3909, n3910, n3912, n3914, 
      n3916, n3917, n3920, n3922, n3923, n3924, n3925, n3926, n3928, n3930, 
      n3932, n3933, n3936, n3938, n3939, n3940, n3941, n3942, n3944, n3946, 
      n3948, n3949, n3952, n3954, n3955, n3956, n3957, n3958, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, 
      n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
      n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, 
      n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, 
      n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
      n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, 
      n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, 
      n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, 
      n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, 
      n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, 
      n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, 
      n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, 
      n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, 
      n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, 
      n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
      n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, 
      n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
      n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, 
      n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
      n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, 
      n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, 
      n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, 
      n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, 
      n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, 
      n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, 
      n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, 
      n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, 
      n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, 
      n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, 
      n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, 
      n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, 
      n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, 
      n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, 
      n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, 
      n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, 
      n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, 
      n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, 
      n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, 
      n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, 
      n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, 
      n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, 
      n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, 
      n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, 
      n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, 
      n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, 
      n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, 
      n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, 
      n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, 
      n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, 
      n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, 
      n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, 
      n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, 
      n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, 
      n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, 
      n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, 
      n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, 
      n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, 
      n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, 
      n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, 
      n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, 
      n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, 
      n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, 
      n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, 
      n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, 
      n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, 
      n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, 
      n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, 
      n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, 
      n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, 
      n9204, n9205, n815, n816, n817, n819, n821, n822, n824, n826, n827, n830,
      n842, n845, n847, n849, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
      n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
      n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
      n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
      n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
      n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
      n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
      n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
      n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
      n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
      n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
      n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
      n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
      n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
      n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
      n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
      n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
      n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
      n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
      n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
      n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
      n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
      n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
      n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
      n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
      n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
      n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
      n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
      n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
      n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
      n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
      n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
      n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
      n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, 
      n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
      n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
      n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
      n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
      n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
      n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
      n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
      n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
      n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
      n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, 
      n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
      n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
      n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, 
      n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
      n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
      n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, 
      n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
      n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
      n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
      n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, 
      n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, 
      n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, 
      n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, 
      n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, 
      n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, 
      n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, 
      n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
      n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, 
      n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, 
      n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, 
      n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, 
      n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
      n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
      n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
      n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, 
      n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, 
      n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, 
      n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, 
      n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, 
      n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, 
      n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, 
      n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, 
      n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, 
      n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, 
      n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, 
      n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
      n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, 
      n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, 
      n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, 
      n2350, n2351, n2352, n2353, n2354, n2355, n9207, n9208, n9209, n9210, 
      n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, 
      n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, 
      n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, 
      n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, 
      n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, 
      n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, 
      n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, 
      n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, 
      n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, 
      n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, 
      n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, 
      n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, 
      n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, 
      n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, 
      n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, 
      n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, 
      n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, 
      n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, 
      n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, 
      n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, 
      n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, 
      n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, 
      n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, 
      n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, 
      n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, 
      n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, 
      n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, 
      n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, 
      n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, 
      n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, 
      n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, 
      n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, 
      n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, 
      n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, 
      n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, 
      n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, 
      n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, 
      n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, 
      n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, 
      n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, 
      n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, 
      n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, 
      n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, 
      n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, 
      n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, 
      n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, 
      n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, 
      n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, 
      n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, 
      n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, 
      n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, 
      n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, 
      n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, 
      n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, 
      n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, 
      n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, 
      n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, 
      n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, 
      n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, 
      n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, 
      n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, 
      n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, 
      n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, 
      n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, 
      n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, 
      n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, 
      n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, 
      n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, 
      n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, 
      n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, 
      n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, 
      n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, 
      n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, 
      n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, 
      n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, 
      n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, 
      n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, 
      n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, 
      n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, 
      n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, 
      n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, 
      n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, 
      n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, 
      n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, 
      n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, 
      n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, 
      n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, 
      n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, 
      n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, 
      n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, 
      n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, 
      n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, 
      n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, 
      n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, 
      n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, 
      n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, 
      n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, 
      n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, 
      n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, 
      n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, 
      n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, 
      n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, 
      n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, 
      n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, 
      n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, 
      n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, 
      n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, 
      n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, 
      n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, 
      n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, 
      n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, 
      n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, 
      n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, 
      n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, 
      n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, 
      n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, 
      n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, 
      n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, 
      n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, 
      n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, 
      n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, 
      n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, 
      n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, 
      n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, 
      n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, 
      n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, 
      n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, 
      n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, 
      n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, 
      n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, 
      n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, 
      n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, 
      n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, 
      n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, 
      n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, 
      n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, 
      n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, 
      n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, 
      n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, 
      n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, 
      n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, 
      n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, 
      n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, 
      n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, 
      n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, 
      n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, 
      n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, 
      n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, 
      n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, 
      n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, 
      n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, 
      n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, 
      n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, 
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, 
      n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, 
      n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, 
      n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, 
      n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, 
      n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, 
      n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350 : 
      std_logic;

begin
   
   U1686 : AND3_X2 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), A3 => RD1, ZN 
                           => n1460);
   U1699 : AND3_X2 port map( A1 => ADD_RD1(3), A2 => n10665, A3 => RD1, ZN => 
                           n1470);
   U1716 : AND3_X2 port map( A1 => ADD_RD1(4), A2 => n10658, A3 => RD1, ZN => 
                           n1458);
   U1722 : AND3_X2 port map( A1 => n10658, A2 => n10665, A3 => RD1, ZN => n1477
                           );
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n3005, CK => CLK, RN => 
                           n9883, Q => n10538, QN => n2102);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n3004, CK => CLK, RN => 
                           n9883, Q => n10539, QN => n2110);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n3003, CK => CLK, RN => 
                           n9883, Q => n10540, QN => n2118);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n3002, CK => CLK, RN => 
                           n9883, Q => n10541, QN => n2126);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n3001, CK => CLK, RN => 
                           n9883, Q => n10542, QN => n2134);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n3000, CK => CLK, RN => 
                           n9883, Q => n10543, QN => n2142);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n2999, CK => CLK, RN => 
                           n9883, Q => n10544, QN => n2150);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n2998, CK => CLK, RN => 
                           n9883, Q => n10545, QN => n2158);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n3133, CK => CLK, RN => 
                           n9883, Q => n10562, QN => n8326);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n3132, CK => CLK, RN => 
                           n9883, Q => n10563, QN => n8325);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n3131, CK => CLK, RN => 
                           n9883, Q => n10564, QN => n8324);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n3130, CK => CLK, RN => 
                           n9883, Q => n10565, QN => n8323);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n3129, CK => CLK, RN => 
                           n9883, Q => n10566, QN => n8322);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n3128, CK => CLK, RN => 
                           n9883, Q => n10567, QN => n8321);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n3127, CK => CLK, RN => 
                           n9883, Q => n10568, QN => n8320);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n3126, CK => CLK, RN => 
                           n9883, Q => n10569, QN => n8319);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n2973, CK => CLK, RN => 
                           n9883, Q => n10554, QN => n8342);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n2972, CK => CLK, RN => 
                           n9883, Q => n10555, QN => n8341);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n2971, CK => CLK, RN => 
                           n9883, Q => n10556, QN => n8340);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n2970, CK => CLK, RN => 
                           n9883, Q => n10557, QN => n8339);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n2969, CK => CLK, RN => 
                           n9883, Q => n10558, QN => n8338);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n2968, CK => CLK, RN => 
                           n9883, Q => n10559, QN => n8337);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n2967, CK => CLK, RN => 
                           n9883, Q => n10560, QN => n8336);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n2966, CK => CLK, RN => 
                           n9883, Q => n10561, QN => n8335);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n3101, CK => CLK, RN => 
                           n9883, Q => n_1063, QN => n8509);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n3100, CK => CLK, RN => 
                           n9883, Q => n_1064, QN => n8508);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n3099, CK => CLK, RN => 
                           n9883, Q => n_1065, QN => n8507);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n3098, CK => CLK, RN => 
                           n9883, Q => n_1066, QN => n8506);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n3097, CK => CLK, RN => 
                           n9883, Q => n_1067, QN => n8505);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n3096, CK => CLK, RN => 
                           n9883, Q => n_1068, QN => n8504);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n3095, CK => CLK, RN => 
                           n9883, Q => n_1069, QN => n8503);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n3094, CK => CLK, RN => 
                           n9883, Q => n_1070, QN => n8502);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n3069, CK => CLK, RN => 
                           n9883, Q => n_1071, QN => n8334);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n3068, CK => CLK, RN => 
                           n9883, Q => n_1072, QN => n8333);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n3067, CK => CLK, RN => 
                           n9883, Q => n_1073, QN => n8332);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n3066, CK => CLK, RN => 
                           n9883, Q => n_1074, QN => n8331);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n3065, CK => CLK, RN => 
                           n9883, Q => n_1075, QN => n8330);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n3064, CK => CLK, RN => 
                           n9883, Q => n_1076, QN => n8329);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n3063, CK => CLK, RN => 
                           n9883, Q => n_1077, QN => n8328);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n3062, CK => CLK, RN => 
                           n9883, Q => n_1078, QN => n8327);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n3165, CK => CLK, RN => 
                           n9883, Q => n_1079, QN => n8597);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n3164, CK => CLK, RN => 
                           n9883, Q => n_1080, QN => n8596);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n3163, CK => CLK, RN => 
                           n9883, Q => n_1081, QN => n8595);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n3162, CK => CLK, RN => 
                           n9883, Q => n_1082, QN => n8594);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n3161, CK => CLK, RN => 
                           n9883, Q => n_1083, QN => n8593);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n3160, CK => CLK, RN => 
                           n9883, Q => n_1084, QN => n8592);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n3159, CK => CLK, RN => 
                           n9883, Q => n_1085, QN => n8591);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n3158, CK => CLK, RN => 
                           n9883, Q => n_1086, QN => n8590);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n3811, CK => CLK, RN => 
                           n9883, Q => n10432, QN => n8448);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n9151, CK => CLK, RN => 
                           n9883, Q => n10280, QN => n2276);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n9023, CK => CLK, RN => 
                           n9883, Q => n10096, QN => n8227);
   REGISTERS_reg_0_9_inst : DFFR_X1 port map( D => n8959, CK => CLK, RN => 
                           n9883, Q => n9944, QN => n2280);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n9102, CK => CLK, RN => 
                           n9883, Q => n10530, QN => n2295);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n9103, CK => CLK, RN => 
                           n9883, Q => n10531, QN => n2303);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n9104, CK => CLK, RN => 
                           n9883, Q => n10532, QN => n2311);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n9105, CK => CLK, RN => 
                           n9883, Q => n10533, QN => n2319);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n9106, CK => CLK, RN => 
                           n9883, Q => n10534, QN => n2327);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n3846, CK => CLK, RN => 
                           n9883, Q => n10498, QN => n8350);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n3862, CK => CLK, RN => 
                           n9883, Q => n10499, QN => n8349);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n3878, CK => CLK, RN => 
                           n9883, Q => n10500, QN => n8348);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n3894, CK => CLK, RN => 
                           n9883, Q => n10501, QN => n8347);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n3910, CK => CLK, RN => 
                           n9883, Q => n10502, QN => n8346);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n3845, CK => CLK, RN => 
                           n9883, Q => n_1087, QN => n8382);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n3861, CK => CLK, RN => 
                           n9883, Q => n_1088, QN => n8381);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n3877, CK => CLK, RN => 
                           n9883, Q => n_1089, QN => n8380);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n3893, CK => CLK, RN => 
                           n9883, Q => n_1090, QN => n8379);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n3909, CK => CLK, RN => 
                           n9883, Q => n_1091, QN => n8378);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n9134, CK => CLK, RN => 
                           n9883, Q => n10626, QN => n8230);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n9135, CK => CLK, RN => 
                           n9883, Q => n10627, QN => n8232);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n9136, CK => CLK, RN => 
                           n9883, Q => n10628, QN => n8234);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n9137, CK => CLK, RN => 
                           n9883, Q => n10629, QN => n8236);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n9138, CK => CLK, RN => 
                           n9883, Q => n10630, QN => n8238);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n3844, CK => CLK, RN => 
                           n9883, Q => n10466, QN => n8414);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n3860, CK => CLK, RN => 
                           n9883, Q => n10467, QN => n8413);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n3876, CK => CLK, RN => 
                           n9883, Q => n10468, QN => n8412);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n3892, CK => CLK, RN => 
                           n9883, Q => n10469, QN => n8411);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n3908, CK => CLK, RN => 
                           n9883, Q => n10470, QN => n8410);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n3459, CK => CLK, RN => 
                           n9883, Q => n10410, QN => n8470);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n3827, CK => CLK, RN => 
                           n9883, Q => n10433, QN => n8447);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n3843, CK => CLK, RN => 
                           n9883, Q => n10434, QN => n8446);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n3859, CK => CLK, RN => 
                           n9883, Q => n10435, QN => n8445);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n3875, CK => CLK, RN => 
                           n9883, Q => n10436, QN => n8444);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n3891, CK => CLK, RN => 
                           n9883, Q => n10437, QN => n8443);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n3907, CK => CLK, RN => 
                           n9883, Q => n10438, QN => n8442);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n3842, CK => CLK, RN => 
                           n9883, Q => n10402, QN => n8517);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n3858, CK => CLK, RN => 
                           n9883, Q => n10403, QN => n8516);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n3874, CK => CLK, RN => 
                           n9883, Q => n10404, QN => n8515);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n3890, CK => CLK, RN => 
                           n9883, Q => n10405, QN => n8514);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n3906, CK => CLK, RN => 
                           n9883, Q => n10406, QN => n8513);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n9173, CK => CLK, RN => 
                           n9883, Q => n10258, QN => n2100);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n9150, CK => CLK, RN => 
                           n9883, Q => n10281, QN => n2284);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n9149, CK => CLK, RN => 
                           n9883, Q => n10282, QN => n2292);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n9148, CK => CLK, RN => 
                           n9883, Q => n10283, QN => n2300);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n9147, CK => CLK, RN => 
                           n9883, Q => n10284, QN => n2308);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n9146, CK => CLK, RN => 
                           n9883, Q => n10285, QN => n2316);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n9145, CK => CLK, RN => 
                           n9883, Q => n10286, QN => n2324);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n9077, CK => CLK, RN => 
                           n9883, Q => n10226, QN => n2107);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n9045, CK => CLK, RN => 
                           n9883, Q => n10074, QN => n8183);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n9022, CK => CLK, RN => 
                           n9883, Q => n10097, QN => n8229);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n9021, CK => CLK, RN => 
                           n9883, Q => n10098, QN => n8231);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n9020, CK => CLK, RN => 
                           n9883, Q => n10099, QN => n8233);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n9019, CK => CLK, RN => 
                           n9883, Q => n10100, QN => n8235);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n9018, CK => CLK, RN => 
                           n9883, Q => n10101, QN => n8237);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n9017, CK => CLK, RN => 
                           n9883, Q => n10102, QN => n8239);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n9013, CK => CLK, RN => 
                           n9883, Q => n10010, QN => n2105);
   REGISTERS_reg_0_31_inst : DFFR_X1 port map( D => n8981, CK => CLK, RN => 
                           n9883, Q => n9922, QN => n2104);
   REGISTERS_reg_0_8_inst : DFFR_X1 port map( D => n8958, CK => CLK, RN => 
                           n9883, Q => n9945, QN => n2288);
   REGISTERS_reg_0_7_inst : DFFR_X1 port map( D => n8957, CK => CLK, RN => 
                           n9883, Q => n9946, QN => n2296);
   REGISTERS_reg_0_6_inst : DFFR_X1 port map( D => n8956, CK => CLK, RN => 
                           n9883, Q => n9947, QN => n2304);
   REGISTERS_reg_0_5_inst : DFFR_X1 port map( D => n8955, CK => CLK, RN => 
                           n9883, Q => n9948, QN => n2312);
   REGISTERS_reg_0_4_inst : DFFR_X1 port map( D => n8954, CK => CLK, RN => 
                           n9883, Q => n9949, QN => n2320);
   REGISTERS_reg_0_3_inst : DFFR_X1 port map( D => n8953, CK => CLK, RN => 
                           n9883, Q => n9950, QN => n2328);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n3840, CK => CLK, RN => 
                           n9883, Q => n10314, QN => n8605);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n3856, CK => CLK, RN => 
                           n9883, Q => n10315, QN => n8604);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n3872, CK => CLK, RN => 
                           n9883, Q => n10316, QN => n8603);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n3888, CK => CLK, RN => 
                           n9883, Q => n10317, QN => n8602);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n3904, CK => CLK, RN => 
                           n9883, Q => n10318, QN => n8601);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n3197, CK => CLK, RN => 
                           n9883, Q => n_1092, QN => n8302);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n3229, CK => CLK, RN => 
                           n9883, Q => n_1093, QN => n8685);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n3837, CK => CLK, RN => 
                           n9883, Q => n10218, QN => n8693);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n3853, CK => CLK, RN => 
                           n9883, Q => n10219, QN => n8692);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n3869, CK => CLK, RN => 
                           n9883, Q => n10220, QN => n8691);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n3885, CK => CLK, RN => 
                           n9883, Q => n10221, QN => n8690);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n3901, CK => CLK, RN => 
                           n9883, Q => n10222, QN => n8689);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n3261, CK => CLK, RN => 
                           n9883, Q => n10578, QN => n8294);
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n3293, CK => CLK, RN => 
                           n9883, Q => n10138, QN => n8773);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n3836, CK => CLK, RN => 
                           n9883, Q => n10130, QN => n2298);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n3852, CK => CLK, RN => 
                           n9883, Q => n10131, QN => n2306);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n3868, CK => CLK, RN => 
                           n9883, Q => n10132, QN => n2314);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n3884, CK => CLK, RN => 
                           n9883, Q => n10133, QN => n2322);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n3900, CK => CLK, RN => 
                           n9883, Q => n10134, QN => n2330);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n3325, CK => CLK, RN => 
                           n9883, Q => n_1094, QN => n8318);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n3357, CK => CLK, RN => 
                           n9883, Q => n_1095, QN => n8829);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n3834, CK => CLK, RN => 
                           n9883, Q => n10066, QN => n8837);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n3850, CK => CLK, RN => 
                           n9883, Q => n10067, QN => n8836);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n3866, CK => CLK, RN => 
                           n9883, Q => n10068, QN => n8835);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n3882, CK => CLK, RN => 
                           n9883, Q => n10069, QN => n8834);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n3898, CK => CLK, RN => 
                           n9883, Q => n10070, QN => n8833);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n3389, CK => CLK, RN => 
                           n9883, Q => n10570, QN => n8310);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n3421, CK => CLK, RN => 
                           n9883, Q => n_1096, QN => n8917);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n3832, CK => CLK, RN => 
                           n9883, Q => n9978, QN => n8925);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n3848, CK => CLK, RN => 
                           n9883, Q => n9979, QN => n8924);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n3864, CK => CLK, RN => 
                           n9883, Q => n9980, QN => n8923);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n3880, CK => CLK, RN => 
                           n9883, Q => n9981, QN => n8922);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n3896, CK => CLK, RN => 
                           n9883, Q => n9982, QN => n8921);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n3175, CK => CLK, RN => 
                           n9883, Q => n_1097, QN => n8639);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n3174, CK => CLK, RN => 
                           n9883, Q => n_1098, QN => n8638);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n3173, CK => CLK, RN => 
                           n9883, Q => n_1099, QN => n8637);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n3172, CK => CLK, RN => 
                           n9883, Q => n_1100, QN => n8636);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n3171, CK => CLK, RN => 
                           n9883, Q => n_1101, QN => n8635);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n3170, CK => CLK, RN => 
                           n9883, Q => n_1102, QN => n8634);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n3169, CK => CLK, RN => 
                           n9883, Q => n_1103, QN => n8633);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n9055, CK => CLK, RN => 
                           n9883, Q => n10248, QN => n2283);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n9054, CK => CLK, RN => 
                           n9883, Q => n10249, QN => n2291);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n9053, CK => CLK, RN => 
                           n9883, Q => n10250, QN => n2299);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n9052, CK => CLK, RN => 
                           n9883, Q => n10251, QN => n2307);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n9051, CK => CLK, RN => 
                           n9883, Q => n10252, QN => n2315);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n9050, CK => CLK, RN => 
                           n9883, Q => n10253, QN => n2323);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n9049, CK => CLK, RN => 
                           n9883, Q => n10254, QN => n2331);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n3303, CK => CLK, RN => 
                           n9883, Q => n_1104, QN => n8783);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n3302, CK => CLK, RN => 
                           n9883, Q => n_1105, QN => n8782);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n3301, CK => CLK, RN => 
                           n9883, Q => n_1106, QN => n8781);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n3300, CK => CLK, RN => 
                           n9883, Q => n_1107, QN => n8780);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n3299, CK => CLK, RN => 
                           n9883, Q => n_1108, QN => n8779);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n3298, CK => CLK, RN => 
                           n9883, Q => n_1109, QN => n8778);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n3297, CK => CLK, RN => 
                           n9883, Q => n_1110, QN => n8777);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n3450, CK => CLK, RN => 
                           n9883, Q => n10042, QN => n8861);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n3802, CK => CLK, RN => 
                           n9883, Q => n10064, QN => n8839);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n3818, CK => CLK, RN => 
                           n9883, Q => n10065, QN => n8838);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n9110, CK => CLK, RN => 
                           n9883, Q => n10546, QN => n8182);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n9132, CK => CLK, RN => 
                           n9883, Q => n10624, QN => n8226);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n9133, CK => CLK, RN => 
                           n9883, Q => n10625, QN => n8228);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n3271, CK => CLK, RN => 
                           n9883, Q => n10160, QN => n8751);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n3270, CK => CLK, RN => 
                           n9883, Q => n10161, QN => n8750);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n3269, CK => CLK, RN => 
                           n9883, Q => n10162, QN => n8749);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n3268, CK => CLK, RN => 
                           n9883, Q => n10163, QN => n8748);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n3267, CK => CLK, RN => 
                           n9883, Q => n10164, QN => n8747);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n3266, CK => CLK, RN => 
                           n9883, Q => n10165, QN => n8746);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n3265, CK => CLK, RN => 
                           n9883, Q => n10166, QN => n8745);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n3399, CK => CLK, RN => 
                           n9883, Q => n_1111, QN => n8895);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n3398, CK => CLK, RN => 
                           n9883, Q => n_1112, QN => n8894);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n3397, CK => CLK, RN => 
                           n9883, Q => n_1113, QN => n8893);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n3396, CK => CLK, RN => 
                           n9883, Q => n_1114, QN => n8892);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n3395, CK => CLK, RN => 
                           n9883, Q => n_1115, QN => n8891);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n3394, CK => CLK, RN => 
                           n9883, Q => n_1116, QN => n8890);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n3393, CK => CLK, RN => 
                           n9883, Q => n_1117, QN => n8889);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n3461, CK => CLK, RN => 
                           n9883, Q => n_1118, QN => n8406);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n3813, CK => CLK, RN => 
                           n9883, Q => n_1119, QN => n8384);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n3829, CK => CLK, RN => 
                           n9883, Q => n_1120, QN => n8383);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n3453, CK => CLK, RN => 
                           n9883, Q => n10194, QN => n8717);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n3805, CK => CLK, RN => 
                           n9883, Q => n10216, QN => n8695);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n3821, CK => CLK, RN => 
                           n9883, Q => n10217, QN => n8694);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n8991, CK => CLK, RN => 
                           n9883, Q => n10032, QN => n2281);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n8990, CK => CLK, RN => 
                           n9883, Q => n10033, QN => n2289);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n8989, CK => CLK, RN => 
                           n9883, Q => n10034, QN => n2297);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n8988, CK => CLK, RN => 
                           n9883, Q => n10035, QN => n2305);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n8987, CK => CLK, RN => 
                           n9883, Q => n10036, QN => n2313);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n8986, CK => CLK, RN => 
                           n9883, Q => n10037, QN => n2321);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n8985, CK => CLK, RN => 
                           n9883, Q => n10038, QN => n2329);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n2997, CK => CLK, RN => 
                           n9883, Q => n10586, QN => n2166);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n2996, CK => CLK, RN => 
                           n9883, Q => n10587, QN => n2174);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n2995, CK => CLK, RN => 
                           n9883, Q => n10588, QN => n2182);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n2994, CK => CLK, RN => 
                           n9883, Q => n10589, QN => n2190);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n2993, CK => CLK, RN => 
                           n9883, Q => n10590, QN => n2198);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n2992, CK => CLK, RN => 
                           n9883, Q => n10591, QN => n2206);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n2991, CK => CLK, RN => 
                           n9883, Q => n10592, QN => n2214);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n2990, CK => CLK, RN => 
                           n9883, Q => n10593, QN => n2222);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n2989, CK => CLK, RN => 
                           n9883, Q => n10594, QN => n2230);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n2988, CK => CLK, RN => 
                           n9883, Q => n10595, QN => n2238);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n2987, CK => CLK, RN => 
                           n9883, Q => n10596, QN => n2246);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n2986, CK => CLK, RN => 
                           n9883, Q => n10597, QN => n2254);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n2985, CK => CLK, RN => 
                           n9883, Q => n10598, QN => n2262);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n2984, CK => CLK, RN => 
                           n9883, Q => n10599, QN => n2270);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n2983, CK => CLK, RN => 
                           n9883, Q => n10600, QN => n2278);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n2982, CK => CLK, RN => 
                           n9883, Q => n10601, QN => n2286);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n2981, CK => CLK, RN => 
                           n9883, Q => n10602, QN => n2294);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n2980, CK => CLK, RN => 
                           n9883, Q => n10603, QN => n2302);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n2979, CK => CLK, RN => 
                           n9883, Q => n10604, QN => n2310);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n2978, CK => CLK, RN => 
                           n9883, Q => n10605, QN => n2318);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n2977, CK => CLK, RN => 
                           n9883, Q => n10606, QN => n2326);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n2976, CK => CLK, RN => 
                           n9883, Q => n10607, QN => n2334);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n2975, CK => CLK, RN => 
                           n9883, Q => n10608, QN => n2342);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n2974, CK => CLK, RN => 
                           n9883, Q => n10609, QN => n2350);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n3460, CK => CLK, RN => 
                           n9883, Q => n10442, QN => n8438);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n3812, CK => CLK, RN => 
                           n9883, Q => n10464, QN => n8416);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n3828, CK => CLK, RN => 
                           n9883, Q => n10465, QN => n8415);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n3125, CK => CLK, RN => 
                           n9883, Q => n10322, QN => n8565);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n3124, CK => CLK, RN => 
                           n9883, Q => n10323, QN => n8564);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n3123, CK => CLK, RN => 
                           n9883, Q => n10324, QN => n8563);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n3122, CK => CLK, RN => 
                           n9883, Q => n10325, QN => n8562);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n3121, CK => CLK, RN => 
                           n9883, Q => n10326, QN => n8561);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n3120, CK => CLK, RN => 
                           n9883, Q => n10327, QN => n8560);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n3119, CK => CLK, RN => 
                           n9883, Q => n10328, QN => n8559);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n3118, CK => CLK, RN => 
                           n9883, Q => n10329, QN => n8558);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n3117, CK => CLK, RN => 
                           n9883, Q => n10330, QN => n8557);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n3116, CK => CLK, RN => 
                           n9883, Q => n10331, QN => n8556);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n3115, CK => CLK, RN => 
                           n9883, Q => n10332, QN => n8555);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n3114, CK => CLK, RN => 
                           n9883, Q => n10333, QN => n8554);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n3113, CK => CLK, RN => 
                           n9883, Q => n10334, QN => n8553);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n3112, CK => CLK, RN => 
                           n9883, Q => n10335, QN => n8552);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n3111, CK => CLK, RN => 
                           n9883, Q => n10336, QN => n8551);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n3110, CK => CLK, RN => 
                           n9883, Q => n10337, QN => n8550);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n3109, CK => CLK, RN => 
                           n9883, Q => n10338, QN => n8549);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n3108, CK => CLK, RN => 
                           n9883, Q => n10339, QN => n8548);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n3107, CK => CLK, RN => 
                           n9883, Q => n10340, QN => n8547);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n3106, CK => CLK, RN => 
                           n9883, Q => n10341, QN => n8546);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n3105, CK => CLK, RN => 
                           n9883, Q => n10342, QN => n8545);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n3104, CK => CLK, RN => 
                           n9883, Q => n10343, QN => n8544);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n3103, CK => CLK, RN => 
                           n9883, Q => n10344, QN => n8543);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n3102, CK => CLK, RN => 
                           n9883, Q => n10345, QN => n8542);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n3456, CK => CLK, RN => 
                           n9883, Q => n10290, QN => n8629);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n3808, CK => CLK, RN => 
                           n9883, Q => n10312, QN => n8607);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n3824, CK => CLK, RN => 
                           n9883, Q => n10313, QN => n8606);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n3239, CK => CLK, RN => 
                           n9883, Q => n10184, QN => n8727);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n3238, CK => CLK, RN => 
                           n9883, Q => n10185, QN => n8726);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n3237, CK => CLK, RN => 
                           n9883, Q => n10186, QN => n8725);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n3236, CK => CLK, RN => 
                           n9883, Q => n10187, QN => n8724);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n3235, CK => CLK, RN => 
                           n9883, Q => n10188, QN => n8723);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n3234, CK => CLK, RN => 
                           n9883, Q => n10189, QN => n8722);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n3233, CK => CLK, RN => 
                           n9883, Q => n10190, QN => n8721);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n3452, CK => CLK, RN => 
                           n9883, Q => n10106, QN => n2106);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n3804, CK => CLK, RN => 
                           n9883, Q => n10128, QN => n2282);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n3820, CK => CLK, RN => 
                           n9883, Q => n10129, QN => n2290);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n3367, CK => CLK, RN => 
                           n9883, Q => n10000, QN => n8871);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n3366, CK => CLK, RN => 
                           n9883, Q => n10001, QN => n8870);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n3365, CK => CLK, RN => 
                           n9883, Q => n10002, QN => n8869);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n3364, CK => CLK, RN => 
                           n9883, Q => n10003, QN => n8868);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n3363, CK => CLK, RN => 
                           n9883, Q => n10004, QN => n8867);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n3362, CK => CLK, RN => 
                           n9883, Q => n10005, QN => n8866);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n3361, CK => CLK, RN => 
                           n9883, Q => n10006, QN => n8865);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n3448, CK => CLK, RN => 
                           n9883, Q => n9954, QN => n8949);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n3800, CK => CLK, RN => 
                           n9883, Q => n9976, QN => n8927);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n3816, CK => CLK, RN => 
                           n9883, Q => n9977, QN => n8926);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n2965, CK => CLK, RN => 
                           n9883, Q => n10634, QN => n8286);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n2964, CK => CLK, RN => 
                           n9883, Q => n10635, QN => n8285);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n2963, CK => CLK, RN => 
                           n9883, Q => n10636, QN => n8284);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n2962, CK => CLK, RN => 
                           n9883, Q => n10637, QN => n8283);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n2961, CK => CLK, RN => 
                           n9883, Q => n10638, QN => n8282);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n2960, CK => CLK, RN => 
                           n9883, Q => n10639, QN => n8281);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n2959, CK => CLK, RN => 
                           n9883, Q => n10640, QN => n8280);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n2958, CK => CLK, RN => 
                           n9883, Q => n10641, QN => n8279);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n2957, CK => CLK, RN => 
                           n9883, Q => n10642, QN => n8278);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n2956, CK => CLK, RN => 
                           n9883, Q => n10643, QN => n8277);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n2955, CK => CLK, RN => 
                           n9883, Q => n10644, QN => n8276);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n2954, CK => CLK, RN => 
                           n9883, Q => n10645, QN => n8275);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n2953, CK => CLK, RN => 
                           n9883, Q => n10646, QN => n8274);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n2952, CK => CLK, RN => 
                           n9883, Q => n10647, QN => n8273);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n2951, CK => CLK, RN => 
                           n9883, Q => n10648, QN => n8272);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n2950, CK => CLK, RN => 
                           n9883, Q => n10649, QN => n8271);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n2949, CK => CLK, RN => 
                           n9883, Q => n10650, QN => n8270);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n2948, CK => CLK, RN => 
                           n9883, Q => n10651, QN => n8269);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n2947, CK => CLK, RN => 
                           n9883, Q => n10652, QN => n8268);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n2946, CK => CLK, RN => 
                           n9883, Q => n10653, QN => n8267);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n2945, CK => CLK, RN => 
                           n9883, Q => n10654, QN => n8266);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n2944, CK => CLK, RN => 
                           n9883, Q => n10655, QN => n8265);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n2943, CK => CLK, RN => 
                           n9883, Q => n10656, QN => n8264);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n2942, CK => CLK, RN => 
                           n9883, Q => n10657, QN => n8263);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n3093, CK => CLK, RN => 
                           n9883, Q => n_1121, QN => n8501);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n3092, CK => CLK, RN => 
                           n9883, Q => n_1122, QN => n8500);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n3091, CK => CLK, RN => 
                           n9883, Q => n_1123, QN => n8499);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n3090, CK => CLK, RN => 
                           n9883, Q => n_1124, QN => n8498);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n3089, CK => CLK, RN => 
                           n9883, Q => n_1125, QN => n8497);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n3088, CK => CLK, RN => 
                           n9883, Q => n_1126, QN => n8496);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n3087, CK => CLK, RN => 
                           n9883, Q => n_1127, QN => n8495);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n3086, CK => CLK, RN => 
                           n9883, Q => n_1128, QN => n8494);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n3085, CK => CLK, RN => 
                           n9883, Q => n_1129, QN => n8493);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n3084, CK => CLK, RN => 
                           n9883, Q => n_1130, QN => n8492);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n3083, CK => CLK, RN => 
                           n9883, Q => n_1131, QN => n8491);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n3082, CK => CLK, RN => 
                           n9883, Q => n_1132, QN => n8490);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n3081, CK => CLK, RN => 
                           n9883, Q => n_1133, QN => n8489);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n3080, CK => CLK, RN => 
                           n9883, Q => n_1134, QN => n8488);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n3079, CK => CLK, RN => 
                           n9883, Q => n_1135, QN => n8487);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n3078, CK => CLK, RN => 
                           n9883, Q => n_1136, QN => n8486);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n3077, CK => CLK, RN => 
                           n9883, Q => n_1137, QN => n8485);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n3076, CK => CLK, RN => 
                           n9883, Q => n_1138, QN => n8484);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n3075, CK => CLK, RN => 
                           n9883, Q => n_1139, QN => n8483);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n3074, CK => CLK, RN => 
                           n9883, Q => n_1140, QN => n8482);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n3073, CK => CLK, RN => 
                           n9883, Q => n_1141, QN => n8481);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n3072, CK => CLK, RN => 
                           n9883, Q => n_1142, QN => n8480);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n3071, CK => CLK, RN => 
                           n9883, Q => n_1143, QN => n8479);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n3070, CK => CLK, RN => 
                           n9883, Q => n_1144, QN => n8478);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n3207, CK => CLK, RN => 
                           n9883, Q => n_1145, QN => n8663);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n3206, CK => CLK, RN => 
                           n9883, Q => n_1146, QN => n8662);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n3205, CK => CLK, RN => 
                           n9883, Q => n_1147, QN => n8661);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n3204, CK => CLK, RN => 
                           n9883, Q => n_1148, QN => n8660);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n3203, CK => CLK, RN => 
                           n9883, Q => n_1149, QN => n8659);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n3202, CK => CLK, RN => 
                           n9883, Q => n_1150, QN => n8658);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n3201, CK => CLK, RN => 
                           n9883, Q => n_1151, QN => n8657);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n3335, CK => CLK, RN => 
                           n9883, Q => n_1152, QN => n8807);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n3334, CK => CLK, RN => 
                           n9883, Q => n_1153, QN => n8806);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n3333, CK => CLK, RN => 
                           n9883, Q => n_1154, QN => n8805);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n3332, CK => CLK, RN => 
                           n9883, Q => n_1155, QN => n8804);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n3331, CK => CLK, RN => 
                           n9883, Q => n_1156, QN => n8803);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n3330, CK => CLK, RN => 
                           n9883, Q => n_1157, QN => n8802);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n3329, CK => CLK, RN => 
                           n9883, Q => n_1158, QN => n8801);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n9078, CK => CLK, RN => 
                           n9883, Q => n10506, QN => n2103);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n9100, CK => CLK, RN => 
                           n9883, Q => n10528, QN => n2279);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n9101, CK => CLK, RN => 
                           n9883, Q => n10529, QN => n2287);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n3061, CK => CLK, RN => 
                           n9883, Q => n_1159, QN => n8262);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n3060, CK => CLK, RN => 
                           n9883, Q => n_1160, QN => n8261);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n3059, CK => CLK, RN => 
                           n9883, Q => n_1161, QN => n8260);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n3058, CK => CLK, RN => 
                           n9883, Q => n_1162, QN => n8259);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n3057, CK => CLK, RN => 
                           n9883, Q => n_1163, QN => n8258);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n3056, CK => CLK, RN => 
                           n9883, Q => n_1164, QN => n8257);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n3055, CK => CLK, RN => 
                           n9883, Q => n_1165, QN => n8256);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n3054, CK => CLK, RN => 
                           n9883, Q => n_1166, QN => n8255);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n3053, CK => CLK, RN => 
                           n9883, Q => n_1167, QN => n8254);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n3052, CK => CLK, RN => 
                           n9883, Q => n_1168, QN => n8253);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n3051, CK => CLK, RN => 
                           n9883, Q => n_1169, QN => n8252);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n3050, CK => CLK, RN => 
                           n9883, Q => n_1170, QN => n8251);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n3049, CK => CLK, RN => 
                           n9883, Q => n_1171, QN => n8250);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n3048, CK => CLK, RN => 
                           n9883, Q => n_1172, QN => n8249);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n3047, CK => CLK, RN => 
                           n9883, Q => n_1173, QN => n8248);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n3046, CK => CLK, RN => 
                           n9883, Q => n_1174, QN => n8247);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n3045, CK => CLK, RN => 
                           n9883, Q => n_1175, QN => n8246);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n3044, CK => CLK, RN => 
                           n9883, Q => n_1176, QN => n8477);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n3043, CK => CLK, RN => 
                           n9883, Q => n_1177, QN => n8476);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n3042, CK => CLK, RN => 
                           n9883, Q => n_1178, QN => n8475);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n3041, CK => CLK, RN => 
                           n9883, Q => n_1179, QN => n8474);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n3040, CK => CLK, RN => 
                           n9883, Q => n_1180, QN => n8473);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n3039, CK => CLK, RN => 
                           n9883, Q => n_1181, QN => n8472);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n3038, CK => CLK, RN => 
                           n9883, Q => n_1182, QN => n8471);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n3462, CK => CLK, RN => 
                           n9883, Q => n10474, QN => n8374);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n3814, CK => CLK, RN => 
                           n9883, Q => n10496, QN => n8352);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n3830, CK => CLK, RN => 
                           n9883, Q => n10497, QN => n8351);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n3458, CK => CLK, RN => 
                           n9883, Q => n10378, QN => n8541);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n3810, CK => CLK, RN => 
                           n9883, Q => n10400, QN => n8519);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n3826, CK => CLK, RN => 
                           n9883, Q => n10401, QN => n8518);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n9205, CK => CLK, RN => 
                           n9878, Q => n10346, QN => n2101);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n3157, CK => CLK, RN => 
                           n9883, Q => n_1183, QN => n8589);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n3156, CK => CLK, RN => 
                           n9883, Q => n_1184, QN => n8588);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n3155, CK => CLK, RN => 
                           n9883, Q => n_1185, QN => n8587);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n3154, CK => CLK, RN => 
                           n9883, Q => n_1186, QN => n8586);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n3153, CK => CLK, RN => 
                           n9883, Q => n_1187, QN => n8585);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n3152, CK => CLK, RN => 
                           n9883, Q => n_1188, QN => n8584);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n3151, CK => CLK, RN => 
                           n9883, Q => n_1189, QN => n8583);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n3150, CK => CLK, RN => 
                           n9883, Q => n_1190, QN => n8582);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n3149, CK => CLK, RN => 
                           n9883, Q => n_1191, QN => n8581);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n3148, CK => CLK, RN => 
                           n9883, Q => n_1192, QN => n8580);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n3147, CK => CLK, RN => 
                           n9883, Q => n_1193, QN => n8579);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n3146, CK => CLK, RN => 
                           n9883, Q => n_1194, QN => n8578);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n3145, CK => CLK, RN => 
                           n9883, Q => n_1195, QN => n8577);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n3144, CK => CLK, RN => 
                           n9883, Q => n_1196, QN => n8576);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n3143, CK => CLK, RN => 
                           n9883, Q => n_1197, QN => n8575);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n3142, CK => CLK, RN => 
                           n9883, Q => n_1198, QN => n8574);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n3141, CK => CLK, RN => 
                           n9883, Q => n_1199, QN => n8573);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n3140, CK => CLK, RN => 
                           n9883, Q => n_1200, QN => n8572);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n3139, CK => CLK, RN => 
                           n9883, Q => n_1201, QN => n8571);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n3138, CK => CLK, RN => 
                           n9883, Q => n_1202, QN => n8570);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n3137, CK => CLK, RN => 
                           n9883, Q => n_1203, QN => n8569);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n3136, CK => CLK, RN => 
                           n9883, Q => n_1204, QN => n8568);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n3135, CK => CLK, RN => 
                           n9883, Q => n_1205, QN => n8567);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n3134, CK => CLK, RN => 
                           n9883, Q => n_1206, QN => n8566);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n9079, CK => CLK, RN => 
                           n9883, Q => n10507, QN => n2111);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n9080, CK => CLK, RN => 
                           n9883, Q => n10508, QN => n2119);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n9081, CK => CLK, RN => 
                           n9883, Q => n10509, QN => n2127);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n9082, CK => CLK, RN => 
                           n9883, Q => n10510, QN => n2135);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n9083, CK => CLK, RN => 
                           n9883, Q => n10511, QN => n2143);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n9084, CK => CLK, RN => 
                           n9883, Q => n10512, QN => n2151);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n9085, CK => CLK, RN => 
                           n9883, Q => n10513, QN => n2159);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n9086, CK => CLK, RN => 
                           n9883, Q => n10514, QN => n2167);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n9087, CK => CLK, RN => 
                           n9883, Q => n10515, QN => n2175);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n9088, CK => CLK, RN => 
                           n9883, Q => n10516, QN => n2183);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n9089, CK => CLK, RN => 
                           n9883, Q => n10517, QN => n2191);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n9090, CK => CLK, RN => 
                           n9883, Q => n10518, QN => n2199);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n9091, CK => CLK, RN => 
                           n9883, Q => n10519, QN => n2207);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n9092, CK => CLK, RN => 
                           n9883, Q => n10520, QN => n2215);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n9093, CK => CLK, RN => 
                           n9883, Q => n10521, QN => n2223);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n9094, CK => CLK, RN => 
                           n9883, Q => n10522, QN => n2231);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n9095, CK => CLK, RN => 
                           n9883, Q => n10523, QN => n2239);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n9096, CK => CLK, RN => 
                           n9883, Q => n10524, QN => n2247);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n9097, CK => CLK, RN => 
                           n9883, Q => n10525, QN => n2255);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n9098, CK => CLK, RN => 
                           n9883, Q => n10526, QN => n2263);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n9099, CK => CLK, RN => 
                           n9883, Q => n10527, QN => n2271);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n9107, CK => CLK, RN => 
                           n9883, Q => n10535, QN => n2335);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n9108, CK => CLK, RN => 
                           n9883, Q => n10536, QN => n2343);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n9109, CK => CLK, RN => 
                           n9883, Q => n10537, QN => n2351);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n3478, CK => CLK, RN => 
                           n9883, Q => n10475, QN => n8373);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n3494, CK => CLK, RN => 
                           n9883, Q => n10476, QN => n8372);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n3510, CK => CLK, RN => 
                           n9883, Q => n10477, QN => n8371);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n3526, CK => CLK, RN => 
                           n9883, Q => n10478, QN => n8370);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n3542, CK => CLK, RN => 
                           n9883, Q => n10479, QN => n8369);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n3558, CK => CLK, RN => 
                           n9883, Q => n10480, QN => n8368);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n3574, CK => CLK, RN => 
                           n9883, Q => n10481, QN => n8367);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n3590, CK => CLK, RN => 
                           n9883, Q => n10482, QN => n8366);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n3606, CK => CLK, RN => 
                           n9883, Q => n10483, QN => n8365);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n3622, CK => CLK, RN => 
                           n9883, Q => n10484, QN => n8364);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n3638, CK => CLK, RN => 
                           n9883, Q => n10485, QN => n8363);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n3654, CK => CLK, RN => 
                           n9883, Q => n10486, QN => n8362);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n3670, CK => CLK, RN => 
                           n9883, Q => n10487, QN => n8361);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n3686, CK => CLK, RN => 
                           n9883, Q => n10488, QN => n8360);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n3702, CK => CLK, RN => 
                           n9883, Q => n10489, QN => n8359);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n3718, CK => CLK, RN => 
                           n9883, Q => n10490, QN => n8358);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n3734, CK => CLK, RN => 
                           n9883, Q => n10491, QN => n8357);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n3750, CK => CLK, RN => 
                           n9883, Q => n10492, QN => n8356);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n3766, CK => CLK, RN => 
                           n9883, Q => n10493, QN => n8355);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n3782, CK => CLK, RN => 
                           n9883, Q => n10494, QN => n8354);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n3798, CK => CLK, RN => 
                           n9883, Q => n10495, QN => n8353);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n3926, CK => CLK, RN => 
                           n9883, Q => n10503, QN => n8345);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n3942, CK => CLK, RN => 
                           n9879, Q => n10504, QN => n8344);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n3958, CK => CLK, RN => 
                           n9883, Q => n10505, QN => n8343);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n3477, CK => CLK, RN => 
                           n9883, Q => n_1207, QN => n8405);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n3493, CK => CLK, RN => 
                           n9883, Q => n_1208, QN => n8404);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n3509, CK => CLK, RN => 
                           n9883, Q => n_1209, QN => n8403);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n3525, CK => CLK, RN => 
                           n9883, Q => n_1210, QN => n8402);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n3541, CK => CLK, RN => 
                           n9883, Q => n_1211, QN => n8401);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n3557, CK => CLK, RN => 
                           n9883, Q => n_1212, QN => n8400);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n3573, CK => CLK, RN => 
                           n9883, Q => n_1213, QN => n8399);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n3589, CK => CLK, RN => 
                           n9883, Q => n_1214, QN => n8398);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n3605, CK => CLK, RN => 
                           n9883, Q => n_1215, QN => n8397);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n3621, CK => CLK, RN => 
                           n9883, Q => n_1216, QN => n8396);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n3637, CK => CLK, RN => 
                           n9883, Q => n_1217, QN => n8395);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n3653, CK => CLK, RN => 
                           n9883, Q => n_1218, QN => n8394);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n3669, CK => CLK, RN => 
                           n9883, Q => n_1219, QN => n8393);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n3685, CK => CLK, RN => 
                           n9883, Q => n_1220, QN => n8392);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n3701, CK => CLK, RN => 
                           n9883, Q => n_1221, QN => n8391);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n3717, CK => CLK, RN => 
                           n9883, Q => n_1222, QN => n8390);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n3733, CK => CLK, RN => 
                           n9883, Q => n_1223, QN => n8389);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n3749, CK => CLK, RN => 
                           n9883, Q => n_1224, QN => n8388);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n3765, CK => CLK, RN => 
                           n9883, Q => n_1225, QN => n8387);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n3781, CK => CLK, RN => 
                           n9883, Q => n_1226, QN => n8386);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n3797, CK => CLK, RN => 
                           n9883, Q => n_1227, QN => n8385);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n3925, CK => CLK, RN => 
                           n9883, Q => n_1228, QN => n8377);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n3941, CK => CLK, RN => 
                           n9879, Q => n_1229, QN => n8376);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n3957, CK => CLK, RN => 
                           n9883, Q => n_1230, QN => n8375);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n9111, CK => CLK, RN => 
                           n9883, Q => n10547, QN => n8184);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n9112, CK => CLK, RN => 
                           n9883, Q => n10548, QN => n8186);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n9113, CK => CLK, RN => 
                           n9883, Q => n10549, QN => n8188);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n9114, CK => CLK, RN => 
                           n9883, Q => n10550, QN => n8190);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n9115, CK => CLK, RN => 
                           n9883, Q => n10551, QN => n8192);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n9116, CK => CLK, RN => 
                           n9883, Q => n10552, QN => n8194);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n9117, CK => CLK, RN => 
                           n9883, Q => n10553, QN => n8196);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n9118, CK => CLK, RN => 
                           n9883, Q => n10610, QN => n8198);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n9119, CK => CLK, RN => 
                           n9883, Q => n10611, QN => n8200);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n9120, CK => CLK, RN => 
                           n9883, Q => n10612, QN => n8202);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n9121, CK => CLK, RN => 
                           n9883, Q => n10613, QN => n8204);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n9122, CK => CLK, RN => 
                           n9883, Q => n10614, QN => n8206);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n9123, CK => CLK, RN => 
                           n9883, Q => n10615, QN => n8208);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n9124, CK => CLK, RN => 
                           n9883, Q => n10616, QN => n8210);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n9125, CK => CLK, RN => 
                           n9883, Q => n10617, QN => n8212);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n9126, CK => CLK, RN => 
                           n9883, Q => n10618, QN => n8214);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n9127, CK => CLK, RN => 
                           n9883, Q => n10619, QN => n8216);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n9128, CK => CLK, RN => 
                           n9883, Q => n10620, QN => n8218);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n9129, CK => CLK, RN => 
                           n9883, Q => n10621, QN => n8220);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n9130, CK => CLK, RN => 
                           n9883, Q => n10622, QN => n8222);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n9131, CK => CLK, RN => 
                           n9883, Q => n10623, QN => n8224);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n9139, CK => CLK, RN => 
                           n9883, Q => n10631, QN => n8240);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n9140, CK => CLK, RN => 
                           n9883, Q => n10632, QN => n8242);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n9141, CK => CLK, RN => 
                           n9883, Q => n10633, QN => n8244);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n3476, CK => CLK, RN => 
                           n9883, Q => n10443, QN => n8437);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n3492, CK => CLK, RN => 
                           n9883, Q => n10444, QN => n8436);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n3508, CK => CLK, RN => 
                           n9883, Q => n10445, QN => n8435);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n3524, CK => CLK, RN => 
                           n9883, Q => n10446, QN => n8434);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n3540, CK => CLK, RN => 
                           n9883, Q => n10447, QN => n8433);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n3556, CK => CLK, RN => 
                           n9883, Q => n10448, QN => n8432);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n3572, CK => CLK, RN => 
                           n9883, Q => n10449, QN => n8431);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n3588, CK => CLK, RN => 
                           n9883, Q => n10450, QN => n8430);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n3604, CK => CLK, RN => 
                           n9883, Q => n10451, QN => n8429);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n3620, CK => CLK, RN => 
                           n9883, Q => n10452, QN => n8428);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n3636, CK => CLK, RN => 
                           n9883, Q => n10453, QN => n8427);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n3652, CK => CLK, RN => 
                           n9883, Q => n10454, QN => n8426);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n3668, CK => CLK, RN => 
                           n9883, Q => n10455, QN => n8425);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n3684, CK => CLK, RN => 
                           n9883, Q => n10456, QN => n8424);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n3700, CK => CLK, RN => 
                           n9883, Q => n10457, QN => n8423);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n3716, CK => CLK, RN => 
                           n9883, Q => n10458, QN => n8422);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n3732, CK => CLK, RN => 
                           n9883, Q => n10459, QN => n8421);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n3748, CK => CLK, RN => 
                           n9883, Q => n10460, QN => n8420);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n3764, CK => CLK, RN => 
                           n9883, Q => n10461, QN => n8419);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n3780, CK => CLK, RN => 
                           n9883, Q => n10462, QN => n8418);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n3796, CK => CLK, RN => 
                           n9883, Q => n10463, QN => n8417);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n3924, CK => CLK, RN => 
                           n9883, Q => n10471, QN => n8409);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n3940, CK => CLK, RN => 
                           n9879, Q => n10472, QN => n8408);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n3956, CK => CLK, RN => 
                           n9883, Q => n10473, QN => n8407);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n3475, CK => CLK, RN => 
                           n9883, Q => n10411, QN => n8469);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n3491, CK => CLK, RN => 
                           n9883, Q => n10412, QN => n8468);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n3507, CK => CLK, RN => 
                           n9883, Q => n10413, QN => n8467);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n3523, CK => CLK, RN => 
                           n9883, Q => n10414, QN => n8466);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n3539, CK => CLK, RN => 
                           n9883, Q => n10415, QN => n8465);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n3555, CK => CLK, RN => 
                           n9883, Q => n10416, QN => n8464);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n3571, CK => CLK, RN => 
                           n9883, Q => n10417, QN => n8463);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n3587, CK => CLK, RN => 
                           n9883, Q => n10418, QN => n8462);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n3603, CK => CLK, RN => 
                           n9883, Q => n10419, QN => n8461);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n3619, CK => CLK, RN => 
                           n9883, Q => n10420, QN => n8460);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n3635, CK => CLK, RN => 
                           n9883, Q => n10421, QN => n8459);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n3651, CK => CLK, RN => 
                           n9883, Q => n10422, QN => n8458);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n3667, CK => CLK, RN => 
                           n9883, Q => n10423, QN => n8457);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n3683, CK => CLK, RN => 
                           n9883, Q => n10424, QN => n8456);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n3699, CK => CLK, RN => 
                           n9883, Q => n10425, QN => n8455);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n3715, CK => CLK, RN => 
                           n9883, Q => n10426, QN => n8454);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n3731, CK => CLK, RN => 
                           n9883, Q => n10427, QN => n8453);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n3747, CK => CLK, RN => 
                           n9883, Q => n10428, QN => n8452);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n3763, CK => CLK, RN => 
                           n9883, Q => n10429, QN => n8451);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n3779, CK => CLK, RN => 
                           n9883, Q => n10430, QN => n8450);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n3795, CK => CLK, RN => 
                           n9883, Q => n10431, QN => n8449);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n3923, CK => CLK, RN => 
                           n9883, Q => n10439, QN => n8441);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n3939, CK => CLK, RN => 
                           n9879, Q => n10440, QN => n8440);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n3955, CK => CLK, RN => 
                           n9883, Q => n10441, QN => n8439);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n3474, CK => CLK, RN => 
                           n9883, Q => n10379, QN => n8540);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n3490, CK => CLK, RN => 
                           n9883, Q => n10380, QN => n8539);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n3506, CK => CLK, RN => 
                           n9883, Q => n10381, QN => n8538);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n3522, CK => CLK, RN => 
                           n9883, Q => n10382, QN => n8537);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n3538, CK => CLK, RN => 
                           n9883, Q => n10383, QN => n8536);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n3554, CK => CLK, RN => 
                           n9883, Q => n10384, QN => n8535);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n3570, CK => CLK, RN => 
                           n9883, Q => n10385, QN => n8534);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n3586, CK => CLK, RN => 
                           n9883, Q => n10386, QN => n8533);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n3602, CK => CLK, RN => 
                           n9883, Q => n10387, QN => n8532);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n3618, CK => CLK, RN => 
                           n9883, Q => n10388, QN => n8531);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n3634, CK => CLK, RN => 
                           n9883, Q => n10389, QN => n8530);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n3650, CK => CLK, RN => 
                           n9883, Q => n10390, QN => n8529);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n3666, CK => CLK, RN => 
                           n9883, Q => n10391, QN => n8528);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n3682, CK => CLK, RN => 
                           n9883, Q => n10392, QN => n8527);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n3698, CK => CLK, RN => 
                           n9883, Q => n10393, QN => n8526);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n3714, CK => CLK, RN => 
                           n9883, Q => n10394, QN => n8525);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n3730, CK => CLK, RN => 
                           n9883, Q => n10395, QN => n8524);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n3746, CK => CLK, RN => 
                           n9883, Q => n10396, QN => n8523);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n3762, CK => CLK, RN => 
                           n9883, Q => n10397, QN => n8522);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n3778, CK => CLK, RN => 
                           n9883, Q => n10398, QN => n8521);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n3794, CK => CLK, RN => 
                           n9883, Q => n10399, QN => n8520);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n3922, CK => CLK, RN => 
                           n9883, Q => n10407, QN => n8512);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n3938, CK => CLK, RN => 
                           n9883, Q => n10408, QN => n8511);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n3954, CK => CLK, RN => 
                           n9883, Q => n10409, QN => n8510);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n9172, CK => CLK, RN => 
                           n9883, Q => n10259, QN => n2108);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n9171, CK => CLK, RN => 
                           n9883, Q => n10260, QN => n2116);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n9170, CK => CLK, RN => 
                           n9883, Q => n10261, QN => n2124);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n9169, CK => CLK, RN => 
                           n9883, Q => n10262, QN => n2132);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n9168, CK => CLK, RN => 
                           n9883, Q => n10263, QN => n2140);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n9167, CK => CLK, RN => 
                           n9883, Q => n10264, QN => n2148);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n9166, CK => CLK, RN => 
                           n9883, Q => n10265, QN => n2156);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n9165, CK => CLK, RN => 
                           n9883, Q => n10266, QN => n2164);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n9164, CK => CLK, RN => 
                           n9883, Q => n10267, QN => n2172);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n9163, CK => CLK, RN => 
                           n9883, Q => n10268, QN => n2180);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n9162, CK => CLK, RN => 
                           n9883, Q => n10269, QN => n2188);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n9161, CK => CLK, RN => 
                           n9883, Q => n10270, QN => n2196);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n9160, CK => CLK, RN => 
                           n9883, Q => n10271, QN => n2204);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n9159, CK => CLK, RN => 
                           n9883, Q => n10272, QN => n2212);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n9158, CK => CLK, RN => 
                           n9883, Q => n10273, QN => n2220);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n9157, CK => CLK, RN => 
                           n9883, Q => n10274, QN => n2228);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n9156, CK => CLK, RN => 
                           n9883, Q => n10275, QN => n2236);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n9155, CK => CLK, RN => 
                           n9883, Q => n10276, QN => n2244);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n9154, CK => CLK, RN => 
                           n9883, Q => n10277, QN => n2252);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n9153, CK => CLK, RN => 
                           n9883, Q => n10278, QN => n2260);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n9152, CK => CLK, RN => 
                           n9883, Q => n10279, QN => n2268);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n9144, CK => CLK, RN => 
                           n9883, Q => n10287, QN => n2332);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n9143, CK => CLK, RN => 
                           n9883, Q => n10288, QN => n2340);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n9142, CK => CLK, RN => 
                           n9883, Q => n10289, QN => n2348);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n9076, CK => CLK, RN => 
                           n9883, Q => n10227, QN => n2115);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n9075, CK => CLK, RN => 
                           n9883, Q => n10228, QN => n2123);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n9074, CK => CLK, RN => 
                           n9883, Q => n10229, QN => n2131);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n9073, CK => CLK, RN => 
                           n9883, Q => n10230, QN => n2139);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n9072, CK => CLK, RN => 
                           n9883, Q => n10231, QN => n2147);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n9071, CK => CLK, RN => 
                           n9883, Q => n10232, QN => n2155);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n9070, CK => CLK, RN => 
                           n9883, Q => n10233, QN => n2163);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n9069, CK => CLK, RN => 
                           n9883, Q => n10234, QN => n2171);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n9068, CK => CLK, RN => 
                           n9883, Q => n10235, QN => n2179);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n9067, CK => CLK, RN => 
                           n9883, Q => n10236, QN => n2187);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n9066, CK => CLK, RN => 
                           n9883, Q => n10237, QN => n2195);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n9065, CK => CLK, RN => 
                           n9883, Q => n10238, QN => n2203);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n9064, CK => CLK, RN => 
                           n9883, Q => n10239, QN => n2211);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n9063, CK => CLK, RN => 
                           n9883, Q => n10240, QN => n2219);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n9062, CK => CLK, RN => 
                           n9883, Q => n10241, QN => n2227);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n9061, CK => CLK, RN => 
                           n9883, Q => n10242, QN => n2235);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n9060, CK => CLK, RN => 
                           n9883, Q => n10243, QN => n2243);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n9059, CK => CLK, RN => 
                           n9883, Q => n10244, QN => n2251);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n9058, CK => CLK, RN => 
                           n9883, Q => n10245, QN => n2259);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n9057, CK => CLK, RN => 
                           n9883, Q => n10246, QN => n2267);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n9056, CK => CLK, RN => 
                           n9883, Q => n10247, QN => n2275);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n9048, CK => CLK, RN => 
                           n9883, Q => n10255, QN => n2339);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n9047, CK => CLK, RN => 
                           n9883, Q => n10256, QN => n2347);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n9046, CK => CLK, RN => 
                           n9883, Q => n10257, QN => n2355);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n9044, CK => CLK, RN => 
                           n9883, Q => n10075, QN => n8185);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n9043, CK => CLK, RN => 
                           n9883, Q => n10076, QN => n8187);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n9042, CK => CLK, RN => 
                           n9883, Q => n10077, QN => n8189);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n9041, CK => CLK, RN => 
                           n9883, Q => n10078, QN => n8191);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n9040, CK => CLK, RN => 
                           n9883, Q => n10079, QN => n8193);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n9039, CK => CLK, RN => 
                           n9883, Q => n10080, QN => n8195);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n9038, CK => CLK, RN => 
                           n9883, Q => n10081, QN => n8197);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n9037, CK => CLK, RN => 
                           n9883, Q => n10082, QN => n8199);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n9036, CK => CLK, RN => 
                           n9883, Q => n10083, QN => n8201);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n9035, CK => CLK, RN => 
                           n9883, Q => n10084, QN => n8203);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n9034, CK => CLK, RN => 
                           n9883, Q => n10085, QN => n8205);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n9033, CK => CLK, RN => 
                           n9883, Q => n10086, QN => n8207);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n9032, CK => CLK, RN => 
                           n9883, Q => n10087, QN => n8209);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n9031, CK => CLK, RN => 
                           n9883, Q => n10088, QN => n8211);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n9030, CK => CLK, RN => 
                           n9883, Q => n10089, QN => n8213);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n9029, CK => CLK, RN => 
                           n9883, Q => n10090, QN => n8215);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n9028, CK => CLK, RN => 
                           n9883, Q => n10091, QN => n8217);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n9027, CK => CLK, RN => 
                           n9883, Q => n10092, QN => n8219);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n9026, CK => CLK, RN => 
                           n9883, Q => n10093, QN => n8221);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n9025, CK => CLK, RN => 
                           n9883, Q => n10094, QN => n8223);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n9024, CK => CLK, RN => 
                           n9883, Q => n10095, QN => n8225);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n9016, CK => CLK, RN => 
                           n9883, Q => n10103, QN => n8241);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n9015, CK => CLK, RN => 
                           n9883, Q => n10104, QN => n8243);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n9014, CK => CLK, RN => 
                           n9883, Q => n10105, QN => n8245);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n9012, CK => CLK, RN => 
                           n9883, Q => n10011, QN => n2113);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n9011, CK => CLK, RN => 
                           n9883, Q => n10012, QN => n2121);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n9010, CK => CLK, RN => 
                           n9883, Q => n10013, QN => n2129);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n9009, CK => CLK, RN => 
                           n9883, Q => n10014, QN => n2137);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n9008, CK => CLK, RN => 
                           n9883, Q => n10015, QN => n2145);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n9007, CK => CLK, RN => 
                           n9883, Q => n10016, QN => n2153);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n9006, CK => CLK, RN => 
                           n9883, Q => n10017, QN => n2161);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n9005, CK => CLK, RN => 
                           n9883, Q => n10018, QN => n2169);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n9004, CK => CLK, RN => 
                           n9883, Q => n10019, QN => n2177);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n9003, CK => CLK, RN => 
                           n9883, Q => n10020, QN => n2185);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n9002, CK => CLK, RN => 
                           n9883, Q => n10021, QN => n2193);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n9001, CK => CLK, RN => 
                           n9883, Q => n10022, QN => n2201);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n9000, CK => CLK, RN => 
                           n9883, Q => n10023, QN => n2209);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n8999, CK => CLK, RN => 
                           n9883, Q => n10024, QN => n2217);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n8998, CK => CLK, RN => 
                           n9883, Q => n10025, QN => n2225);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n8997, CK => CLK, RN => 
                           n9883, Q => n10026, QN => n2233);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n8996, CK => CLK, RN => 
                           n9883, Q => n10027, QN => n2241);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n8995, CK => CLK, RN => 
                           n9883, Q => n10028, QN => n2249);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n8994, CK => CLK, RN => 
                           n9883, Q => n10029, QN => n2257);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n8993, CK => CLK, RN => 
                           n9883, Q => n10030, QN => n2265);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n8992, CK => CLK, RN => 
                           n9883, Q => n10031, QN => n2273);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n8984, CK => CLK, RN => 
                           n9883, Q => n10039, QN => n2337);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n8983, CK => CLK, RN => 
                           n9883, Q => n10040, QN => n2345);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n8982, CK => CLK, RN => 
                           n9883, Q => n10041, QN => n2353);
   REGISTERS_reg_0_30_inst : DFFR_X1 port map( D => n8980, CK => CLK, RN => 
                           n9883, Q => n9923, QN => n2112);
   REGISTERS_reg_0_29_inst : DFFR_X1 port map( D => n8979, CK => CLK, RN => 
                           n9883, Q => n9924, QN => n2120);
   REGISTERS_reg_0_28_inst : DFFR_X1 port map( D => n8978, CK => CLK, RN => 
                           n9883, Q => n9925, QN => n2128);
   REGISTERS_reg_0_27_inst : DFFR_X1 port map( D => n8977, CK => CLK, RN => 
                           n9883, Q => n9926, QN => n2136);
   REGISTERS_reg_0_26_inst : DFFR_X1 port map( D => n8976, CK => CLK, RN => 
                           n9883, Q => n9927, QN => n2144);
   REGISTERS_reg_0_25_inst : DFFR_X1 port map( D => n8975, CK => CLK, RN => 
                           n9883, Q => n9928, QN => n2152);
   REGISTERS_reg_0_24_inst : DFFR_X1 port map( D => n8974, CK => CLK, RN => 
                           n9883, Q => n9929, QN => n2160);
   REGISTERS_reg_0_23_inst : DFFR_X1 port map( D => n8973, CK => CLK, RN => 
                           n9883, Q => n9930, QN => n2168);
   REGISTERS_reg_0_22_inst : DFFR_X1 port map( D => n8972, CK => CLK, RN => 
                           n9883, Q => n9931, QN => n2176);
   REGISTERS_reg_0_21_inst : DFFR_X1 port map( D => n8971, CK => CLK, RN => 
                           n9883, Q => n9932, QN => n2184);
   REGISTERS_reg_0_20_inst : DFFR_X1 port map( D => n8970, CK => CLK, RN => 
                           n9883, Q => n9933, QN => n2192);
   REGISTERS_reg_0_19_inst : DFFR_X1 port map( D => n8969, CK => CLK, RN => 
                           n9883, Q => n9934, QN => n2200);
   REGISTERS_reg_0_18_inst : DFFR_X1 port map( D => n8968, CK => CLK, RN => 
                           n9883, Q => n9935, QN => n2208);
   REGISTERS_reg_0_17_inst : DFFR_X1 port map( D => n8967, CK => CLK, RN => 
                           n9883, Q => n9936, QN => n2216);
   REGISTERS_reg_0_16_inst : DFFR_X1 port map( D => n8966, CK => CLK, RN => 
                           n9883, Q => n9937, QN => n2224);
   REGISTERS_reg_0_15_inst : DFFR_X1 port map( D => n8965, CK => CLK, RN => 
                           n9883, Q => n9938, QN => n2232);
   REGISTERS_reg_0_14_inst : DFFR_X1 port map( D => n8964, CK => CLK, RN => 
                           n9883, Q => n9939, QN => n2240);
   REGISTERS_reg_0_13_inst : DFFR_X1 port map( D => n8963, CK => CLK, RN => 
                           n9883, Q => n9940, QN => n2248);
   REGISTERS_reg_0_12_inst : DFFR_X1 port map( D => n8962, CK => CLK, RN => 
                           n9883, Q => n9941, QN => n2256);
   REGISTERS_reg_0_11_inst : DFFR_X1 port map( D => n8961, CK => CLK, RN => 
                           n9883, Q => n9942, QN => n2264);
   REGISTERS_reg_0_10_inst : DFFR_X1 port map( D => n8960, CK => CLK, RN => 
                           n9883, Q => n9943, QN => n2272);
   REGISTERS_reg_0_2_inst : DFFR_X1 port map( D => n8952, CK => CLK, RN => 
                           n9883, Q => n9951, QN => n2336);
   REGISTERS_reg_0_1_inst : DFFR_X1 port map( D => n8951, CK => CLK, RN => 
                           n9883, Q => n9952, QN => n2344);
   REGISTERS_reg_0_0_inst : DFFR_X1 port map( D => n8950, CK => CLK, RN => 
                           n9883, Q => n9953, QN => n2352);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n3472, CK => CLK, RN => 
                           n9883, Q => n10291, QN => n8628);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n3488, CK => CLK, RN => 
                           n9883, Q => n10292, QN => n8627);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n3504, CK => CLK, RN => 
                           n9883, Q => n10293, QN => n8626);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n3520, CK => CLK, RN => 
                           n9883, Q => n10294, QN => n8625);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n3536, CK => CLK, RN => 
                           n9883, Q => n10295, QN => n8624);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n3552, CK => CLK, RN => 
                           n9883, Q => n10296, QN => n8623);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n3568, CK => CLK, RN => 
                           n9883, Q => n10297, QN => n8622);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n3584, CK => CLK, RN => 
                           n9883, Q => n10298, QN => n8621);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n3600, CK => CLK, RN => 
                           n9883, Q => n10299, QN => n8620);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n3616, CK => CLK, RN => 
                           n9883, Q => n10300, QN => n8619);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n3632, CK => CLK, RN => 
                           n9883, Q => n10301, QN => n8618);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n3648, CK => CLK, RN => 
                           n9883, Q => n10302, QN => n8617);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n3664, CK => CLK, RN => 
                           n9883, Q => n10303, QN => n8616);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n3680, CK => CLK, RN => 
                           n9883, Q => n10304, QN => n8615);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n3696, CK => CLK, RN => 
                           n9883, Q => n10305, QN => n8614);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n3712, CK => CLK, RN => 
                           n9883, Q => n10306, QN => n8613);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n3728, CK => CLK, RN => 
                           n9883, Q => n10307, QN => n8612);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n3744, CK => CLK, RN => 
                           n9883, Q => n10308, QN => n8611);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n3760, CK => CLK, RN => 
                           n9883, Q => n10309, QN => n8610);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n3776, CK => CLK, RN => 
                           n9883, Q => n10310, QN => n8609);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n3792, CK => CLK, RN => 
                           n9883, Q => n10311, QN => n8608);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n3920, CK => CLK, RN => 
                           n9883, Q => n10319, QN => n8600);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n3936, CK => CLK, RN => 
                           n9883, Q => n10320, QN => n8599);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n3952, CK => CLK, RN => 
                           n9883, Q => n10321, QN => n8598);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n3196, CK => CLK, RN => 
                           n9883, Q => n_1231, QN => n8301);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n3195, CK => CLK, RN => 
                           n9883, Q => n_1232, QN => n8300);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n3194, CK => CLK, RN => 
                           n9883, Q => n_1233, QN => n8299);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n3193, CK => CLK, RN => 
                           n9883, Q => n_1234, QN => n8298);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n3192, CK => CLK, RN => 
                           n9883, Q => n_1235, QN => n8297);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n3191, CK => CLK, RN => 
                           n9883, Q => n_1236, QN => n8296);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n3190, CK => CLK, RN => 
                           n9883, Q => n_1237, QN => n8295);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n3189, CK => CLK, RN => 
                           n9883, Q => n_1238, QN => n8653);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n3188, CK => CLK, RN => 
                           n9883, Q => n_1239, QN => n8652);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n3187, CK => CLK, RN => 
                           n9883, Q => n_1240, QN => n8651);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n3186, CK => CLK, RN => 
                           n9883, Q => n_1241, QN => n8650);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n3185, CK => CLK, RN => 
                           n9883, Q => n_1242, QN => n8649);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n3184, CK => CLK, RN => 
                           n9883, Q => n_1243, QN => n8648);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n3183, CK => CLK, RN => 
                           n9883, Q => n_1244, QN => n8647);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n3182, CK => CLK, RN => 
                           n9883, Q => n_1245, QN => n8646);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n3181, CK => CLK, RN => 
                           n9883, Q => n_1246, QN => n8645);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n3180, CK => CLK, RN => 
                           n9883, Q => n_1247, QN => n8644);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n3179, CK => CLK, RN => 
                           n9883, Q => n_1248, QN => n8643);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n3178, CK => CLK, RN => 
                           n9883, Q => n_1249, QN => n8642);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n3177, CK => CLK, RN => 
                           n9883, Q => n_1250, QN => n8641);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n3176, CK => CLK, RN => 
                           n9883, Q => n_1251, QN => n8640);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n3168, CK => CLK, RN => 
                           n9883, Q => n_1252, QN => n8632);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n3167, CK => CLK, RN => 
                           n9883, Q => n_1253, QN => n8631);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n3166, CK => CLK, RN => 
                           n9883, Q => n_1254, QN => n8630);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n3228, CK => CLK, RN => 
                           n9883, Q => n_1255, QN => n8684);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n3227, CK => CLK, RN => 
                           n9883, Q => n_1256, QN => n8683);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n3226, CK => CLK, RN => 
                           n9883, Q => n_1257, QN => n8682);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n3225, CK => CLK, RN => 
                           n9883, Q => n_1258, QN => n8681);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n3224, CK => CLK, RN => 
                           n9883, Q => n_1259, QN => n8680);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n3223, CK => CLK, RN => 
                           n9883, Q => n_1260, QN => n8679);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n3222, CK => CLK, RN => 
                           n9883, Q => n_1261, QN => n8678);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n3221, CK => CLK, RN => 
                           n9883, Q => n_1262, QN => n8677);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n3220, CK => CLK, RN => 
                           n9883, Q => n_1263, QN => n8676);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n3219, CK => CLK, RN => 
                           n9883, Q => n_1264, QN => n8675);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n3218, CK => CLK, RN => 
                           n9883, Q => n_1265, QN => n8674);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n3217, CK => CLK, RN => 
                           n9883, Q => n_1266, QN => n8673);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n3216, CK => CLK, RN => 
                           n9883, Q => n_1267, QN => n8672);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n3215, CK => CLK, RN => 
                           n9883, Q => n_1268, QN => n8671);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n3214, CK => CLK, RN => 
                           n9883, Q => n_1269, QN => n8670);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n3213, CK => CLK, RN => 
                           n9883, Q => n_1270, QN => n8669);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n3212, CK => CLK, RN => 
                           n9883, Q => n_1271, QN => n8668);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n3211, CK => CLK, RN => 
                           n9883, Q => n_1272, QN => n8667);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n3210, CK => CLK, RN => 
                           n9883, Q => n_1273, QN => n8666);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n3209, CK => CLK, RN => 
                           n9883, Q => n_1274, QN => n8665);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n3208, CK => CLK, RN => 
                           n9883, Q => n_1275, QN => n8664);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n3200, CK => CLK, RN => 
                           n9883, Q => n_1276, QN => n8656);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n3199, CK => CLK, RN => 
                           n9883, Q => n_1277, QN => n8655);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n3198, CK => CLK, RN => 
                           n9883, Q => n_1278, QN => n8654);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n3469, CK => CLK, RN => 
                           n9883, Q => n10195, QN => n8716);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n3485, CK => CLK, RN => 
                           n9883, Q => n10196, QN => n8715);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n3501, CK => CLK, RN => 
                           n9883, Q => n10197, QN => n8714);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n3517, CK => CLK, RN => 
                           n9883, Q => n10198, QN => n8713);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n3533, CK => CLK, RN => 
                           n9883, Q => n10199, QN => n8712);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n3549, CK => CLK, RN => 
                           n9883, Q => n10200, QN => n8711);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n3565, CK => CLK, RN => 
                           n9883, Q => n10201, QN => n8710);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n3581, CK => CLK, RN => 
                           n9883, Q => n10202, QN => n8709);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n3597, CK => CLK, RN => 
                           n9883, Q => n10203, QN => n8708);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n3613, CK => CLK, RN => 
                           n9883, Q => n10204, QN => n8707);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n3629, CK => CLK, RN => 
                           n9883, Q => n10205, QN => n8706);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n3645, CK => CLK, RN => 
                           n9883, Q => n10206, QN => n8705);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n3661, CK => CLK, RN => 
                           n9883, Q => n10207, QN => n8704);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n3677, CK => CLK, RN => 
                           n9883, Q => n10208, QN => n8703);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n3693, CK => CLK, RN => 
                           n9883, Q => n10209, QN => n8702);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n3709, CK => CLK, RN => 
                           n9883, Q => n10210, QN => n8701);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n3725, CK => CLK, RN => 
                           n9883, Q => n10211, QN => n8700);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n3741, CK => CLK, RN => 
                           n9883, Q => n10212, QN => n8699);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n3757, CK => CLK, RN => 
                           n9883, Q => n10213, QN => n8698);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n3773, CK => CLK, RN => 
                           n9883, Q => n10214, QN => n8697);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n3789, CK => CLK, RN => 
                           n9883, Q => n10215, QN => n8696);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n3917, CK => CLK, RN => 
                           n9883, Q => n10223, QN => n8688);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n3933, CK => CLK, RN => 
                           n9883, Q => n10224, QN => n8687);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n3949, CK => CLK, RN => 
                           n9883, Q => n10225, QN => n8686);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n3260, CK => CLK, RN => 
                           n9883, Q => n10579, QN => n8293);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n3259, CK => CLK, RN => 
                           n9883, Q => n10580, QN => n8292);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n3258, CK => CLK, RN => 
                           n9883, Q => n10581, QN => n8291);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n3257, CK => CLK, RN => 
                           n9883, Q => n10582, QN => n8290);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n3256, CK => CLK, RN => 
                           n9883, Q => n10583, QN => n8289);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n3255, CK => CLK, RN => 
                           n9883, Q => n10584, QN => n8288);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n3254, CK => CLK, RN => 
                           n9883, Q => n10585, QN => n8287);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n3253, CK => CLK, RN => 
                           n9883, Q => n10170, QN => n8741);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n3252, CK => CLK, RN => 
                           n9883, Q => n10171, QN => n8740);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n3251, CK => CLK, RN => 
                           n9883, Q => n10172, QN => n8739);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n3250, CK => CLK, RN => 
                           n9883, Q => n10173, QN => n8738);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n3249, CK => CLK, RN => 
                           n9883, Q => n10174, QN => n8737);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n3248, CK => CLK, RN => 
                           n9883, Q => n10175, QN => n8736);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n3247, CK => CLK, RN => 
                           n9883, Q => n10176, QN => n8735);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n3246, CK => CLK, RN => 
                           n9883, Q => n10177, QN => n8734);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n3245, CK => CLK, RN => 
                           n9883, Q => n10178, QN => n8733);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n3244, CK => CLK, RN => 
                           n9883, Q => n10179, QN => n8732);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n3243, CK => CLK, RN => 
                           n9883, Q => n10180, QN => n8731);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n3242, CK => CLK, RN => 
                           n9883, Q => n10181, QN => n8730);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n3241, CK => CLK, RN => 
                           n9883, Q => n10182, QN => n8729);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n3240, CK => CLK, RN => 
                           n9883, Q => n10183, QN => n8728);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n3232, CK => CLK, RN => 
                           n9883, Q => n10191, QN => n8720);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n3231, CK => CLK, RN => 
                           n9883, Q => n10192, QN => n8719);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n3230, CK => CLK, RN => 
                           n9883, Q => n10193, QN => n8718);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n3292, CK => CLK, RN => 
                           n9883, Q => n10139, QN => n8772);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n3291, CK => CLK, RN => 
                           n9883, Q => n10140, QN => n8771);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n3290, CK => CLK, RN => 
                           n9883, Q => n10141, QN => n8770);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n3289, CK => CLK, RN => 
                           n9883, Q => n10142, QN => n8769);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n3288, CK => CLK, RN => 
                           n9883, Q => n10143, QN => n8768);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n3287, CK => CLK, RN => 
                           n9883, Q => n10144, QN => n8767);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n3286, CK => CLK, RN => 
                           n9883, Q => n10145, QN => n8766);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n3285, CK => CLK, RN => 
                           n9883, Q => n10146, QN => n8765);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n3284, CK => CLK, RN => 
                           n9883, Q => n10147, QN => n8764);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n3283, CK => CLK, RN => 
                           n9883, Q => n10148, QN => n8763);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n3282, CK => CLK, RN => 
                           n9883, Q => n10149, QN => n8762);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n3281, CK => CLK, RN => 
                           n9883, Q => n10150, QN => n8761);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n3280, CK => CLK, RN => 
                           n9883, Q => n10151, QN => n8760);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n3279, CK => CLK, RN => 
                           n9883, Q => n10152, QN => n8759);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n3278, CK => CLK, RN => 
                           n9883, Q => n10153, QN => n8758);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n3277, CK => CLK, RN => 
                           n9883, Q => n10154, QN => n8757);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n3276, CK => CLK, RN => 
                           n9883, Q => n10155, QN => n8756);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n3275, CK => CLK, RN => 
                           n9883, Q => n10156, QN => n8755);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n3274, CK => CLK, RN => 
                           n9883, Q => n10157, QN => n8754);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n3273, CK => CLK, RN => 
                           n9883, Q => n10158, QN => n8753);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n3272, CK => CLK, RN => 
                           n9883, Q => n10159, QN => n8752);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n3264, CK => CLK, RN => 
                           n9883, Q => n10167, QN => n8744);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n3263, CK => CLK, RN => 
                           n9883, Q => n10168, QN => n8743);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n3262, CK => CLK, RN => 
                           n9883, Q => n10169, QN => n8742);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n3468, CK => CLK, RN => 
                           n9883, Q => n10107, QN => n2114);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n3484, CK => CLK, RN => 
                           n9883, Q => n10108, QN => n2122);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n3500, CK => CLK, RN => 
                           n9883, Q => n10109, QN => n2130);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n3516, CK => CLK, RN => 
                           n9883, Q => n10110, QN => n2138);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n3532, CK => CLK, RN => 
                           n9883, Q => n10111, QN => n2146);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n3548, CK => CLK, RN => 
                           n9883, Q => n10112, QN => n2154);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n3564, CK => CLK, RN => 
                           n9883, Q => n10113, QN => n2162);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n3580, CK => CLK, RN => 
                           n9883, Q => n10114, QN => n2170);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n3596, CK => CLK, RN => 
                           n9883, Q => n10115, QN => n2178);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n3612, CK => CLK, RN => 
                           n9883, Q => n10116, QN => n2186);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n3628, CK => CLK, RN => 
                           n9883, Q => n10117, QN => n2194);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n3644, CK => CLK, RN => 
                           n9883, Q => n10118, QN => n2202);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n3660, CK => CLK, RN => 
                           n9883, Q => n10119, QN => n2210);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n3676, CK => CLK, RN => 
                           n9883, Q => n10120, QN => n2218);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n3692, CK => CLK, RN => 
                           n9883, Q => n10121, QN => n2226);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n3708, CK => CLK, RN => 
                           n9883, Q => n10122, QN => n2234);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n3724, CK => CLK, RN => 
                           n9883, Q => n10123, QN => n2242);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n3740, CK => CLK, RN => 
                           n9883, Q => n10124, QN => n2250);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n3756, CK => CLK, RN => 
                           n9883, Q => n10125, QN => n2258);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n3772, CK => CLK, RN => 
                           n9883, Q => n10126, QN => n2266);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n3788, CK => CLK, RN => 
                           n9883, Q => n10127, QN => n2274);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n3916, CK => CLK, RN => 
                           n9883, Q => n10135, QN => n2338);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n3932, CK => CLK, RN => 
                           n9883, Q => n10136, QN => n2346);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n3948, CK => CLK, RN => 
                           n9883, Q => n10137, QN => n2354);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n3324, CK => CLK, RN => 
                           n9883, Q => n_1279, QN => n8317);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n3323, CK => CLK, RN => 
                           n9883, Q => n_1280, QN => n8316);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n3322, CK => CLK, RN => 
                           n9883, Q => n_1281, QN => n8315);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n3321, CK => CLK, RN => 
                           n9883, Q => n_1282, QN => n8314);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n3320, CK => CLK, RN => 
                           n9883, Q => n_1283, QN => n8313);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n3319, CK => CLK, RN => 
                           n9883, Q => n_1284, QN => n8312);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n3318, CK => CLK, RN => 
                           n9883, Q => n_1285, QN => n8311);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n3317, CK => CLK, RN => 
                           n9883, Q => n_1286, QN => n8797);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n3316, CK => CLK, RN => 
                           n9883, Q => n_1287, QN => n8796);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n3315, CK => CLK, RN => 
                           n9883, Q => n_1288, QN => n8795);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n3314, CK => CLK, RN => 
                           n9883, Q => n_1289, QN => n8794);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n3313, CK => CLK, RN => 
                           n9883, Q => n_1290, QN => n8793);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n3312, CK => CLK, RN => 
                           n9883, Q => n_1291, QN => n8792);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n3311, CK => CLK, RN => 
                           n9883, Q => n_1292, QN => n8791);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n3310, CK => CLK, RN => 
                           n9883, Q => n_1293, QN => n8790);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n3309, CK => CLK, RN => 
                           n9883, Q => n_1294, QN => n8789);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n3308, CK => CLK, RN => 
                           n9883, Q => n_1295, QN => n8788);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n3307, CK => CLK, RN => 
                           n9883, Q => n_1296, QN => n8787);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n3306, CK => CLK, RN => 
                           n9883, Q => n_1297, QN => n8786);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n3305, CK => CLK, RN => 
                           n9883, Q => n_1298, QN => n8785);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n3304, CK => CLK, RN => 
                           n9883, Q => n_1299, QN => n8784);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n3296, CK => CLK, RN => 
                           n9883, Q => n_1300, QN => n8776);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n3295, CK => CLK, RN => 
                           n9883, Q => n_1301, QN => n8775);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n3294, CK => CLK, RN => 
                           n9883, Q => n_1302, QN => n8774);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n3356, CK => CLK, RN => 
                           n9883, Q => n_1303, QN => n8828);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n3355, CK => CLK, RN => 
                           n9883, Q => n_1304, QN => n8827);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n3354, CK => CLK, RN => 
                           n9883, Q => n_1305, QN => n8826);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n3353, CK => CLK, RN => 
                           n9883, Q => n_1306, QN => n8825);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n3352, CK => CLK, RN => 
                           n9883, Q => n_1307, QN => n8824);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n3351, CK => CLK, RN => 
                           n9883, Q => n_1308, QN => n8823);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n3350, CK => CLK, RN => 
                           n9883, Q => n_1309, QN => n8822);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n3349, CK => CLK, RN => 
                           n9883, Q => n_1310, QN => n8821);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n3348, CK => CLK, RN => 
                           n9883, Q => n_1311, QN => n8820);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n3347, CK => CLK, RN => 
                           n9883, Q => n_1312, QN => n8819);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n3346, CK => CLK, RN => 
                           n9883, Q => n_1313, QN => n8818);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n3345, CK => CLK, RN => 
                           n9883, Q => n_1314, QN => n8817);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n3344, CK => CLK, RN => 
                           n9883, Q => n_1315, QN => n8816);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n3343, CK => CLK, RN => 
                           n9883, Q => n_1316, QN => n8815);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n3342, CK => CLK, RN => 
                           n9883, Q => n_1317, QN => n8814);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n3341, CK => CLK, RN => 
                           n9883, Q => n_1318, QN => n8813);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n3340, CK => CLK, RN => 
                           n9883, Q => n_1319, QN => n8812);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n3339, CK => CLK, RN => 
                           n9883, Q => n_1320, QN => n8811);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n3338, CK => CLK, RN => 
                           n9883, Q => n_1321, QN => n8810);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n3337, CK => CLK, RN => 
                           n9883, Q => n_1322, QN => n8809);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n3336, CK => CLK, RN => 
                           n9883, Q => n_1323, QN => n8808);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n3328, CK => CLK, RN => 
                           n9883, Q => n_1324, QN => n8800);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n3327, CK => CLK, RN => 
                           n9883, Q => n_1325, QN => n8799);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n3326, CK => CLK, RN => 
                           n9883, Q => n_1326, QN => n8798);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n3466, CK => CLK, RN => 
                           n9883, Q => n10043, QN => n8860);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n3482, CK => CLK, RN => 
                           n9883, Q => n10044, QN => n8859);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n3498, CK => CLK, RN => 
                           n9883, Q => n10045, QN => n8858);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n3514, CK => CLK, RN => 
                           n9883, Q => n10046, QN => n8857);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n3530, CK => CLK, RN => 
                           n9883, Q => n10047, QN => n8856);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n3546, CK => CLK, RN => 
                           n9883, Q => n10048, QN => n8855);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n3562, CK => CLK, RN => 
                           n9883, Q => n10049, QN => n8854);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n3578, CK => CLK, RN => 
                           n9883, Q => n10050, QN => n8853);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n3594, CK => CLK, RN => 
                           n9883, Q => n10051, QN => n8852);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n3610, CK => CLK, RN => 
                           n9883, Q => n10052, QN => n8851);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n3626, CK => CLK, RN => 
                           n9883, Q => n10053, QN => n8850);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n3642, CK => CLK, RN => 
                           n9883, Q => n10054, QN => n8849);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n3658, CK => CLK, RN => 
                           n9883, Q => n10055, QN => n8848);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n3674, CK => CLK, RN => 
                           n9883, Q => n10056, QN => n8847);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n3690, CK => CLK, RN => 
                           n9883, Q => n10057, QN => n8846);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n3706, CK => CLK, RN => 
                           n9883, Q => n10058, QN => n8845);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n3722, CK => CLK, RN => 
                           n9883, Q => n10059, QN => n8844);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n3738, CK => CLK, RN => 
                           n9883, Q => n10060, QN => n8843);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n3754, CK => CLK, RN => 
                           n9883, Q => n10061, QN => n8842);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n3770, CK => CLK, RN => 
                           n9883, Q => n10062, QN => n8841);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n3786, CK => CLK, RN => 
                           n9883, Q => n10063, QN => n8840);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n3914, CK => CLK, RN => 
                           n9883, Q => n10071, QN => n8832);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n3930, CK => CLK, RN => 
                           n9883, Q => n10072, QN => n8831);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n3946, CK => CLK, RN => 
                           n9883, Q => n10073, QN => n8830);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n3388, CK => CLK, RN => 
                           n9883, Q => n10571, QN => n8309);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n3387, CK => CLK, RN => 
                           n9883, Q => n10572, QN => n8308);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n3386, CK => CLK, RN => 
                           n9883, Q => n10573, QN => n8307);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n3385, CK => CLK, RN => 
                           n9883, Q => n10574, QN => n8306);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n3384, CK => CLK, RN => 
                           n9883, Q => n10575, QN => n8305);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n3383, CK => CLK, RN => 
                           n9883, Q => n10576, QN => n8304);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n3382, CK => CLK, RN => 
                           n9883, Q => n10577, QN => n8303);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n3381, CK => CLK, RN => 
                           n9883, Q => n9986, QN => n8885);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n3380, CK => CLK, RN => 
                           n9883, Q => n9987, QN => n8884);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n3379, CK => CLK, RN => 
                           n9883, Q => n9988, QN => n8883);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n3378, CK => CLK, RN => 
                           n9883, Q => n9989, QN => n8882);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n3377, CK => CLK, RN => 
                           n9883, Q => n9990, QN => n8881);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n3376, CK => CLK, RN => 
                           n9883, Q => n9991, QN => n8880);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n3375, CK => CLK, RN => 
                           n9883, Q => n9992, QN => n8879);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n3374, CK => CLK, RN => 
                           n9883, Q => n9993, QN => n8878);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n3373, CK => CLK, RN => 
                           n9883, Q => n9994, QN => n8877);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n3372, CK => CLK, RN => 
                           n9883, Q => n9995, QN => n8876);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n3371, CK => CLK, RN => 
                           n9883, Q => n9996, QN => n8875);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n3370, CK => CLK, RN => 
                           n9883, Q => n9997, QN => n8874);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n3369, CK => CLK, RN => 
                           n9883, Q => n9998, QN => n8873);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n3368, CK => CLK, RN => 
                           n9883, Q => n9999, QN => n8872);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n3360, CK => CLK, RN => 
                           n9883, Q => n10007, QN => n8864);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n3359, CK => CLK, RN => 
                           n9883, Q => n10008, QN => n8863);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n3358, CK => CLK, RN => 
                           n9883, Q => n10009, QN => n8862);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n3420, CK => CLK, RN => 
                           n9883, Q => n_1327, QN => n8916);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n3419, CK => CLK, RN => 
                           n9883, Q => n_1328, QN => n8915);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n3418, CK => CLK, RN => 
                           n9883, Q => n_1329, QN => n8914);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n3417, CK => CLK, RN => 
                           n9883, Q => n_1330, QN => n8913);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n3416, CK => CLK, RN => 
                           n9883, Q => n_1331, QN => n8912);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n3415, CK => CLK, RN => 
                           n9883, Q => n_1332, QN => n8911);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n3414, CK => CLK, RN => 
                           n9883, Q => n_1333, QN => n8910);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n3413, CK => CLK, RN => 
                           n9883, Q => n_1334, QN => n8909);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n3412, CK => CLK, RN => 
                           n9883, Q => n_1335, QN => n8908);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n3411, CK => CLK, RN => 
                           n9883, Q => n_1336, QN => n8907);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n3410, CK => CLK, RN => 
                           n9883, Q => n_1337, QN => n8906);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n3409, CK => CLK, RN => 
                           n9883, Q => n_1338, QN => n8905);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n3408, CK => CLK, RN => 
                           n9883, Q => n_1339, QN => n8904);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n3407, CK => CLK, RN => 
                           n9883, Q => n_1340, QN => n8903);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n3406, CK => CLK, RN => 
                           n9883, Q => n_1341, QN => n8902);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n3405, CK => CLK, RN => 
                           n9883, Q => n_1342, QN => n8901);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n3404, CK => CLK, RN => 
                           n9883, Q => n_1343, QN => n8900);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n3403, CK => CLK, RN => 
                           n9883, Q => n_1344, QN => n8899);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n3402, CK => CLK, RN => 
                           n9883, Q => n_1345, QN => n8898);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n3401, CK => CLK, RN => 
                           n9883, Q => n_1346, QN => n8897);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n3400, CK => CLK, RN => 
                           n9883, Q => n_1347, QN => n8896);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n3392, CK => CLK, RN => 
                           n9883, Q => n_1348, QN => n8888);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n3391, CK => CLK, RN => 
                           n9883, Q => n_1349, QN => n8887);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n3390, CK => CLK, RN => 
                           n9883, Q => n_1350, QN => n8886);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n3464, CK => CLK, RN => 
                           n9883, Q => n9955, QN => n8948);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n3480, CK => CLK, RN => 
                           n9883, Q => n9956, QN => n8947);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n3496, CK => CLK, RN => 
                           n9883, Q => n9957, QN => n8946);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n3512, CK => CLK, RN => 
                           n9883, Q => n9958, QN => n8945);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n3528, CK => CLK, RN => 
                           n9883, Q => n9959, QN => n8944);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n3544, CK => CLK, RN => 
                           n9883, Q => n9960, QN => n8943);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n3560, CK => CLK, RN => 
                           n9883, Q => n9961, QN => n8942);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n3576, CK => CLK, RN => 
                           n9883, Q => n9962, QN => n8941);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n3592, CK => CLK, RN => 
                           n9883, Q => n9963, QN => n8940);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n3608, CK => CLK, RN => 
                           n9883, Q => n9964, QN => n8939);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n3624, CK => CLK, RN => 
                           n9883, Q => n9965, QN => n8938);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n3640, CK => CLK, RN => 
                           n9883, Q => n9966, QN => n8937);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n3656, CK => CLK, RN => 
                           n9883, Q => n9967, QN => n8936);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n3672, CK => CLK, RN => 
                           n9883, Q => n9968, QN => n8935);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n3688, CK => CLK, RN => 
                           n9883, Q => n9969, QN => n8934);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n3704, CK => CLK, RN => 
                           n9883, Q => n9970, QN => n8933);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n3720, CK => CLK, RN => 
                           n9883, Q => n9971, QN => n8932);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n3736, CK => CLK, RN => 
                           n9883, Q => n9972, QN => n8931);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n3752, CK => CLK, RN => 
                           n9883, Q => n9973, QN => n8930);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n3768, CK => CLK, RN => 
                           n9883, Q => n9974, QN => n8929);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n3784, CK => CLK, RN => 
                           n9883, Q => n9975, QN => n8928);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n3912, CK => CLK, RN => 
                           n9883, Q => n9983, QN => n8920);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n3928, CK => CLK, RN => 
                           n9883, Q => n9984, QN => n8919);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n3944, CK => CLK, RN => 
                           n9883, Q => n9985, QN => n8918);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n9204, CK => CLK, RN => 
                           n9878, Q => n10347, QN => n2109);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n9203, CK => CLK, RN => 
                           n9878, Q => n10348, QN => n2117);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n9202, CK => CLK, RN => 
                           n9878, Q => n10349, QN => n2125);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n9201, CK => CLK, RN => 
                           n9878, Q => n10350, QN => n2133);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n9200, CK => CLK, RN => 
                           n9883, Q => n10351, QN => n2141);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n9199, CK => CLK, RN => 
                           n9878, Q => n10352, QN => n2149);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n9198, CK => CLK, RN => 
                           n9878, Q => n10353, QN => n2157);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n9183, CK => CLK, RN => 
                           n9883, Q => n10368, QN => n2277);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n9197, CK => CLK, RN => 
                           n9877, Q => n10354, QN => n2165);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n9196, CK => CLK, RN => 
                           n9877, Q => n10355, QN => n2173);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n9195, CK => CLK, RN => 
                           n9877, Q => n10356, QN => n2181);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n9194, CK => CLK, RN => 
                           n9877, Q => n10357, QN => n2189);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n9193, CK => CLK, RN => 
                           n9883, Q => n10358, QN => n2197);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n9192, CK => CLK, RN => 
                           n9883, Q => n10359, QN => n2205);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n9191, CK => CLK, RN => 
                           n9883, Q => n10360, QN => n2213);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n9190, CK => CLK, RN => 
                           n9877, Q => n10361, QN => n2221);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n9189, CK => CLK, RN => 
                           n9877, Q => n10362, QN => n2229);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n9188, CK => CLK, RN => 
                           n9883, Q => n10363, QN => n2237);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n9187, CK => CLK, RN => 
                           n9883, Q => n10364, QN => n2245);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n9186, CK => CLK, RN => 
                           n9883, Q => n10365, QN => n2253);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n9185, CK => CLK, RN => 
                           n9882, Q => n10366, QN => n2261);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n9184, CK => CLK, RN => 
                           n9883, Q => n10367, QN => n2269);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n9182, CK => CLK, RN => 
                           n9883, Q => n10369, QN => n2285);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n9181, CK => CLK, RN => 
                           n9883, Q => n10370, QN => n2293);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n9180, CK => CLK, RN => 
                           n9883, Q => n10371, QN => n2301);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n9179, CK => CLK, RN => 
                           n9883, Q => n10372, QN => n2309);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n9178, CK => CLK, RN => 
                           n9883, Q => n10373, QN => n2317);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n9177, CK => CLK, RN => 
                           n9877, Q => n10374, QN => n2325);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n9176, CK => CLK, RN => 
                           n9883, Q => n10375, QN => n2333);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n9175, CK => CLK, RN => 
                           n9883, Q => n10376, QN => n2341);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n9174, CK => CLK, RN => 
                           n9877, Q => n10377, QN => n2349);
   U2 : AND2_X1 port map( A1 => n822, A2 => n816, ZN => n9207);
   U3 : AND2_X1 port map( A1 => n819, A2 => n816, ZN => n9208);
   U4 : AND2_X1 port map( A1 => n824, A2 => n821, ZN => n9209);
   U5 : AND2_X1 port map( A1 => n827, A2 => n816, ZN => n9210);
   U6 : AND2_X1 port map( A1 => n824, A2 => n816, ZN => n9211);
   U7 : AND2_X1 port map( A1 => n827, A2 => n821, ZN => n9212);
   U8 : AND2_X1 port map( A1 => n847, A2 => n826, ZN => n9213);
   U9 : AND2_X1 port map( A1 => n842, A2 => n816, ZN => n9214);
   U10 : AND2_X1 port map( A1 => n842, A2 => n830, ZN => n9215);
   U11 : AND2_X1 port map( A1 => n847, A2 => n816, ZN => n9216);
   U12 : AND2_X1 port map( A1 => n847, A2 => n830, ZN => n9217);
   U13 : AND2_X1 port map( A1 => n842, A2 => n821, ZN => n9218);
   U14 : AND2_X1 port map( A1 => n845, A2 => n816, ZN => n9219);
   U15 : AND2_X1 port map( A1 => n845, A2 => n826, ZN => n9220);
   U16 : AND2_X1 port map( A1 => n845, A2 => n830, ZN => n9221);
   U17 : AND2_X1 port map( A1 => n847, A2 => n821, ZN => n9222);
   U18 : AND2_X1 port map( A1 => n845, A2 => n821, ZN => n9223);
   U19 : AND2_X1 port map( A1 => n842, A2 => n826, ZN => n9224);
   U20 : AND2_X1 port map( A1 => n821, A2 => n819, ZN => n9225);
   U21 : AND2_X1 port map( A1 => n826, A2 => n822, ZN => n9226);
   U22 : AND2_X1 port map( A1 => n830, A2 => n827, ZN => n9227);
   U23 : AND2_X1 port map( A1 => n821, A2 => n817, ZN => n9228);
   U24 : AND2_X1 port map( A1 => n830, A2 => n824, ZN => n9229);
   U25 : AND2_X1 port map( A1 => n830, A2 => n822, ZN => n9230);
   U26 : AND2_X1 port map( A1 => n821, A2 => n822, ZN => n9231);
   U27 : AND2_X1 port map( A1 => n826, A2 => n819, ZN => n9232);
   U28 : AND2_X1 port map( A1 => n826, A2 => n824, ZN => n9233);
   U29 : AND2_X1 port map( A1 => n826, A2 => n827, ZN => n9234);
   U30 : AND2_X1 port map( A1 => n826, A2 => n817, ZN => n9235);
   U31 : AND2_X1 port map( A1 => n830, A2 => n817, ZN => n9236);
   U32 : AND2_X1 port map( A1 => n830, A2 => n819, ZN => n9237);
   U33 : INV_X32 port map( A => n9876, ZN => n9883);
   U34 : CLKBUF_X1 port map( A => RESET, Z => n9876);
   U35 : INV_X1 port map( A => n9646, ZN => n9636);
   U36 : INV_X1 port map( A => n9646, ZN => n9637);
   U37 : INV_X1 port map( A => n9558, ZN => n9549);
   U38 : INV_X1 port map( A => n9536, ZN => n9526);
   U39 : INV_X1 port map( A => n9536, ZN => n9527);
   U40 : INV_X1 port map( A => n9855, ZN => n9846);
   U41 : INV_X1 port map( A => n9547, ZN => n9537);
   U42 : INV_X1 port map( A => n9547, ZN => n9538);
   U43 : INV_X1 port map( A => n9855, ZN => n9845);
   U44 : INV_X1 port map( A => n9844, ZN => n9835);
   U45 : INV_X1 port map( A => n9844, ZN => n9834);
   U46 : INV_X1 port map( A => n9789, ZN => n9780);
   U47 : INV_X1 port map( A => n9789, ZN => n9779);
   U48 : INV_X1 port map( A => n9778, ZN => n9769);
   U49 : INV_X1 port map( A => n9778, ZN => n9768);
   U50 : INV_X1 port map( A => n9767, ZN => n9758);
   U51 : INV_X1 port map( A => n9767, ZN => n9757);
   U52 : INV_X1 port map( A => n9756, ZN => n9747);
   U53 : INV_X1 port map( A => n9756, ZN => n9746);
   U54 : INV_X1 port map( A => n9558, ZN => n9548);
   U55 : INV_X1 port map( A => n9569, ZN => n9559);
   U56 : INV_X1 port map( A => n9569, ZN => n9560);
   U57 : INV_X1 port map( A => n9745, ZN => n9736);
   U58 : INV_X1 port map( A => n9745, ZN => n9735);
   U59 : INV_X1 port map( A => n9580, ZN => n9570);
   U60 : INV_X1 port map( A => n9580, ZN => n9571);
   U61 : INV_X1 port map( A => n9591, ZN => n9581);
   U62 : INV_X1 port map( A => n9591, ZN => n9582);
   U63 : INV_X1 port map( A => n9734, ZN => n9725);
   U64 : INV_X1 port map( A => n9734, ZN => n9724);
   U65 : INV_X1 port map( A => n9866, ZN => n9856);
   U66 : INV_X1 port map( A => n9866, ZN => n9857);
   U67 : INV_X1 port map( A => n9602, ZN => n9592);
   U68 : INV_X1 port map( A => n9602, ZN => n9593);
   U69 : INV_X1 port map( A => n9613, ZN => n9603);
   U70 : INV_X1 port map( A => n9613, ZN => n9604);
   U71 : INV_X1 port map( A => n9833, ZN => n9823);
   U72 : INV_X1 port map( A => n9833, ZN => n9824);
   U73 : INV_X1 port map( A => n9723, ZN => n9714);
   U74 : INV_X1 port map( A => n9723, ZN => n9713);
   U75 : INV_X1 port map( A => n9624, ZN => n9614);
   U76 : INV_X1 port map( A => n9624, ZN => n9615);
   U77 : INV_X1 port map( A => n9635, ZN => n9625);
   U78 : INV_X1 port map( A => n9635, ZN => n9626);
   U79 : INV_X1 port map( A => n9712, ZN => n9703);
   U80 : INV_X1 port map( A => n9712, ZN => n9702);
   U81 : INV_X1 port map( A => n9822, ZN => n9812);
   U82 : INV_X1 port map( A => n9822, ZN => n9813);
   U83 : INV_X1 port map( A => n9657, ZN => n9647);
   U84 : INV_X1 port map( A => n9657, ZN => n9648);
   U85 : INV_X1 port map( A => n9701, ZN => n9692);
   U86 : INV_X1 port map( A => n9701, ZN => n9691);
   U87 : INV_X1 port map( A => n9811, ZN => n9801);
   U88 : INV_X1 port map( A => n9811, ZN => n9802);
   U89 : INV_X1 port map( A => n9668, ZN => n9658);
   U90 : INV_X1 port map( A => n9668, ZN => n9659);
   U91 : INV_X1 port map( A => n9679, ZN => n9669);
   U92 : INV_X1 port map( A => n9679, ZN => n9670);
   U93 : INV_X1 port map( A => n9690, ZN => n9681);
   U94 : INV_X1 port map( A => n9690, ZN => n9680);
   U95 : INV_X1 port map( A => n9800, ZN => n9790);
   U96 : INV_X1 port map( A => n9800, ZN => n9791);
   U97 : BUF_X1 port map( A => n9229, Z => n9646);
   U98 : BUF_X1 port map( A => n9229, Z => n9639);
   U99 : BUF_X1 port map( A => n9229, Z => n9638);
   U100 : BUF_X1 port map( A => n9643, Z => n9645);
   U101 : BUF_X1 port map( A => n9642, Z => n9644);
   U102 : BUF_X1 port map( A => n9229, Z => n9643);
   U103 : BUF_X1 port map( A => n9229, Z => n9642);
   U104 : BUF_X1 port map( A => n9229, Z => n9641);
   U105 : BUF_X1 port map( A => n9229, Z => n9640);
   U106 : INV_X1 port map( A => n9875, ZN => n9867);
   U107 : INV_X1 port map( A => n9875, ZN => n9868);
   U108 : BUF_X1 port map( A => n9210, Z => n9745);
   U109 : BUF_X1 port map( A => n9207, Z => n9591);
   U110 : BUF_X1 port map( A => n9208, Z => n9866);
   U111 : BUF_X1 port map( A => n9222, Z => n9536);
   U112 : BUF_X1 port map( A => n9223, Z => n9547);
   U113 : BUF_X1 port map( A => n9209, Z => n9844);
   U114 : BUF_X1 port map( A => n9212, Z => n9789);
   U115 : BUF_X1 port map( A => n9218, Z => n9767);
   U116 : BUF_X1 port map( A => n9211, Z => n9558);
   U117 : BUF_X1 port map( A => n9216, Z => n9569);
   U118 : BUF_X1 port map( A => n9219, Z => n9580);
   U119 : BUF_X1 port map( A => n9214, Z => n9734);
   U120 : BUF_X1 port map( A => n9213, Z => n9613);
   U121 : BUF_X1 port map( A => n9220, Z => n9624);
   U122 : BUF_X1 port map( A => n9224, Z => n9712);
   U123 : BUF_X1 port map( A => n9217, Z => n9657);
   U124 : BUF_X1 port map( A => n9221, Z => n9668);
   U125 : BUF_X1 port map( A => n9215, Z => n9690);
   U126 : BUF_X1 port map( A => n9231, Z => n9855);
   U127 : BUF_X1 port map( A => n9228, Z => n9778);
   U128 : BUF_X1 port map( A => n9225, Z => n9756);
   U129 : BUF_X1 port map( A => n9233, Z => n9602);
   U130 : BUF_X1 port map( A => n9234, Z => n9833);
   U131 : BUF_X1 port map( A => n9235, Z => n9723);
   U132 : BUF_X1 port map( A => n9226, Z => n9635);
   U133 : BUF_X1 port map( A => n9232, Z => n9822);
   U134 : BUF_X1 port map( A => n9227, Z => n9701);
   U135 : BUF_X1 port map( A => n9236, Z => n9811);
   U136 : BUF_X1 port map( A => n9230, Z => n9679);
   U137 : BUF_X1 port map( A => n9237, Z => n9800);
   U138 : BUF_X1 port map( A => n9211, Z => n9555);
   U139 : BUF_X1 port map( A => n9211, Z => n9554);
   U140 : BUF_X1 port map( A => n9211, Z => n9553);
   U141 : BUF_X1 port map( A => n9211, Z => n9552);
   U142 : BUF_X1 port map( A => n9209, Z => n9838);
   U143 : BUF_X1 port map( A => n9209, Z => n9840);
   U144 : BUF_X1 port map( A => n9840, Z => n9842);
   U145 : BUF_X1 port map( A => n9839, Z => n9843);
   U146 : BUF_X1 port map( A => n9212, Z => n9783);
   U147 : BUF_X1 port map( A => n9212, Z => n9784);
   U148 : BUF_X1 port map( A => n9212, Z => n9785);
   U149 : BUF_X1 port map( A => n9212, Z => n9786);
   U150 : BUF_X1 port map( A => n9784, Z => n9787);
   U151 : BUF_X1 port map( A => n9785, Z => n9788);
   U152 : BUF_X1 port map( A => n9210, Z => n9742);
   U153 : BUF_X1 port map( A => n9585, Z => n9589);
   U154 : BUF_X1 port map( A => n9207, Z => n9588);
   U155 : BUF_X1 port map( A => n9207, Z => n9587);
   U156 : BUF_X1 port map( A => n9207, Z => n9586);
   U157 : BUF_X1 port map( A => n9207, Z => n9585);
   U158 : BUF_X1 port map( A => n9207, Z => n9584);
   U159 : BUF_X1 port map( A => n9207, Z => n9583);
   U160 : BUF_X1 port map( A => n9860, Z => n9865);
   U161 : BUF_X1 port map( A => n9859, Z => n9864);
   U162 : BUF_X1 port map( A => n9208, Z => n9863);
   U163 : BUF_X1 port map( A => n9208, Z => n9862);
   U164 : BUF_X1 port map( A => n9208, Z => n9861);
   U165 : BUF_X1 port map( A => n9208, Z => n9860);
   U166 : BUF_X1 port map( A => n9208, Z => n9859);
   U167 : BUF_X1 port map( A => n9208, Z => n9858);
   U168 : BUF_X1 port map( A => n9530, Z => n9535);
   U169 : BUF_X1 port map( A => n9533, Z => n9534);
   U170 : BUF_X1 port map( A => n9222, Z => n9533);
   U171 : BUF_X1 port map( A => n9222, Z => n9532);
   U172 : BUF_X1 port map( A => n9222, Z => n9531);
   U173 : BUF_X1 port map( A => n9222, Z => n9530);
   U174 : BUF_X1 port map( A => n9541, Z => n9546);
   U175 : BUF_X1 port map( A => n9544, Z => n9545);
   U176 : BUF_X1 port map( A => n9223, Z => n9544);
   U177 : BUF_X1 port map( A => n9223, Z => n9543);
   U178 : BUF_X1 port map( A => n9223, Z => n9542);
   U179 : BUF_X1 port map( A => n9223, Z => n9541);
   U180 : BUF_X1 port map( A => n9220, Z => n9617);
   U181 : BUF_X1 port map( A => n9220, Z => n9616);
   U182 : BUF_X1 port map( A => n9221, Z => n9661);
   U183 : BUF_X1 port map( A => n9221, Z => n9660);
   U184 : BUF_X1 port map( A => n9219, Z => n9573);
   U185 : BUF_X1 port map( A => n9219, Z => n9572);
   U186 : BUF_X1 port map( A => n9211, Z => n9551);
   U187 : BUF_X1 port map( A => n9211, Z => n9550);
   U188 : BUF_X1 port map( A => n9222, Z => n9529);
   U189 : BUF_X1 port map( A => n9222, Z => n9528);
   U190 : BUF_X1 port map( A => n9223, Z => n9540);
   U191 : BUF_X1 port map( A => n9223, Z => n9539);
   U192 : BUF_X1 port map( A => n9209, Z => n9836);
   U193 : BUF_X1 port map( A => n9209, Z => n9837);
   U194 : BUF_X1 port map( A => n9209, Z => n9839);
   U195 : BUF_X1 port map( A => n9209, Z => n9841);
   U196 : BUF_X1 port map( A => n9212, Z => n9781);
   U197 : BUF_X1 port map( A => n9212, Z => n9782);
   U198 : BUF_X1 port map( A => n9218, Z => n9759);
   U199 : BUF_X1 port map( A => n9218, Z => n9760);
   U200 : BUF_X1 port map( A => n9218, Z => n9761);
   U201 : BUF_X1 port map( A => n9218, Z => n9762);
   U202 : BUF_X1 port map( A => n9218, Z => n9763);
   U203 : BUF_X1 port map( A => n9218, Z => n9764);
   U204 : BUF_X1 port map( A => n9762, Z => n9765);
   U205 : BUF_X1 port map( A => n9763, Z => n9766);
   U206 : BUF_X1 port map( A => n9552, Z => n9557);
   U207 : BUF_X1 port map( A => n9555, Z => n9556);
   U208 : BUF_X1 port map( A => n9563, Z => n9568);
   U209 : BUF_X1 port map( A => n9566, Z => n9567);
   U210 : BUF_X1 port map( A => n9216, Z => n9566);
   U211 : BUF_X1 port map( A => n9216, Z => n9565);
   U212 : BUF_X1 port map( A => n9216, Z => n9564);
   U213 : BUF_X1 port map( A => n9216, Z => n9563);
   U214 : BUF_X1 port map( A => n9216, Z => n9562);
   U215 : BUF_X1 port map( A => n9216, Z => n9561);
   U216 : BUF_X1 port map( A => n9210, Z => n9737);
   U217 : BUF_X1 port map( A => n9210, Z => n9738);
   U218 : BUF_X1 port map( A => n9210, Z => n9739);
   U219 : BUF_X1 port map( A => n9210, Z => n9740);
   U220 : BUF_X1 port map( A => n9210, Z => n9741);
   U221 : BUF_X1 port map( A => n9742, Z => n9743);
   U222 : BUF_X1 port map( A => n9740, Z => n9744);
   U223 : BUF_X1 port map( A => n9588, Z => n9590);
   U224 : BUF_X1 port map( A => n9574, Z => n9579);
   U225 : BUF_X1 port map( A => n9577, Z => n9578);
   U226 : BUF_X1 port map( A => n9219, Z => n9577);
   U227 : BUF_X1 port map( A => n9219, Z => n9576);
   U228 : BUF_X1 port map( A => n9219, Z => n9575);
   U229 : BUF_X1 port map( A => n9219, Z => n9574);
   U230 : BUF_X1 port map( A => n9214, Z => n9726);
   U231 : BUF_X1 port map( A => n9214, Z => n9727);
   U232 : BUF_X1 port map( A => n9214, Z => n9728);
   U233 : BUF_X1 port map( A => n9214, Z => n9729);
   U234 : BUF_X1 port map( A => n9214, Z => n9730);
   U235 : BUF_X1 port map( A => n9214, Z => n9731);
   U236 : BUF_X1 port map( A => n9726, Z => n9732);
   U237 : BUF_X1 port map( A => n9727, Z => n9733);
   U238 : BUF_X1 port map( A => n9610, Z => n9612);
   U239 : BUF_X1 port map( A => n9609, Z => n9611);
   U240 : BUF_X1 port map( A => n9213, Z => n9610);
   U241 : BUF_X1 port map( A => n9213, Z => n9609);
   U242 : BUF_X1 port map( A => n9213, Z => n9608);
   U243 : BUF_X1 port map( A => n9213, Z => n9607);
   U244 : BUF_X1 port map( A => n9213, Z => n9606);
   U245 : BUF_X1 port map( A => n9213, Z => n9605);
   U246 : BUF_X1 port map( A => n9617, Z => n9623);
   U247 : BUF_X1 port map( A => n9616, Z => n9622);
   U248 : BUF_X1 port map( A => n9220, Z => n9621);
   U249 : BUF_X1 port map( A => n9220, Z => n9620);
   U250 : BUF_X1 port map( A => n9220, Z => n9619);
   U251 : BUF_X1 port map( A => n9220, Z => n9618);
   U252 : BUF_X1 port map( A => n9224, Z => n9704);
   U253 : BUF_X1 port map( A => n9224, Z => n9705);
   U254 : BUF_X1 port map( A => n9224, Z => n9706);
   U255 : BUF_X1 port map( A => n9224, Z => n9707);
   U256 : BUF_X1 port map( A => n9224, Z => n9708);
   U257 : BUF_X1 port map( A => n9224, Z => n9709);
   U258 : BUF_X1 port map( A => n9707, Z => n9710);
   U259 : BUF_X1 port map( A => n9708, Z => n9711);
   U260 : BUF_X1 port map( A => n9651, Z => n9656);
   U261 : BUF_X1 port map( A => n9650, Z => n9655);
   U262 : BUF_X1 port map( A => n9217, Z => n9654);
   U263 : BUF_X1 port map( A => n9217, Z => n9653);
   U264 : BUF_X1 port map( A => n9217, Z => n9652);
   U265 : BUF_X1 port map( A => n9217, Z => n9651);
   U266 : BUF_X1 port map( A => n9217, Z => n9650);
   U267 : BUF_X1 port map( A => n9217, Z => n9649);
   U268 : BUF_X1 port map( A => n9661, Z => n9667);
   U269 : BUF_X1 port map( A => n9660, Z => n9666);
   U270 : BUF_X1 port map( A => n9221, Z => n9665);
   U271 : BUF_X1 port map( A => n9221, Z => n9664);
   U272 : BUF_X1 port map( A => n9221, Z => n9663);
   U273 : BUF_X1 port map( A => n9221, Z => n9662);
   U274 : BUF_X1 port map( A => n9215, Z => n9682);
   U275 : BUF_X1 port map( A => n9215, Z => n9683);
   U276 : BUF_X1 port map( A => n9215, Z => n9684);
   U277 : BUF_X1 port map( A => n9215, Z => n9685);
   U278 : BUF_X1 port map( A => n9215, Z => n9686);
   U279 : BUF_X1 port map( A => n9215, Z => n9687);
   U280 : BUF_X1 port map( A => n9685, Z => n9688);
   U281 : BUF_X1 port map( A => n9686, Z => n9689);
   U282 : BUF_X1 port map( A => n9231, Z => n9847);
   U283 : BUF_X1 port map( A => n9231, Z => n9848);
   U284 : BUF_X1 port map( A => n9231, Z => n9849);
   U285 : BUF_X1 port map( A => n9231, Z => n9850);
   U286 : BUF_X1 port map( A => n9231, Z => n9851);
   U287 : BUF_X1 port map( A => n9231, Z => n9852);
   U288 : BUF_X1 port map( A => n9233, Z => n9595);
   U289 : BUF_X1 port map( A => n9233, Z => n9594);
   U290 : BUF_X1 port map( A => n9850, Z => n9853);
   U291 : BUF_X1 port map( A => n9851, Z => n9854);
   U292 : BUF_X1 port map( A => n9228, Z => n9770);
   U293 : BUF_X1 port map( A => n9228, Z => n9771);
   U294 : BUF_X1 port map( A => n9228, Z => n9772);
   U295 : BUF_X1 port map( A => n9228, Z => n9773);
   U296 : BUF_X1 port map( A => n9228, Z => n9774);
   U297 : BUF_X1 port map( A => n9228, Z => n9775);
   U298 : BUF_X1 port map( A => n9773, Z => n9776);
   U299 : BUF_X1 port map( A => n9774, Z => n9777);
   U300 : BUF_X1 port map( A => n9225, Z => n9748);
   U301 : BUF_X1 port map( A => n9225, Z => n9749);
   U302 : BUF_X1 port map( A => n9225, Z => n9750);
   U303 : BUF_X1 port map( A => n9225, Z => n9751);
   U304 : BUF_X1 port map( A => n9225, Z => n9752);
   U305 : BUF_X1 port map( A => n9225, Z => n9753);
   U306 : BUF_X1 port map( A => n9751, Z => n9754);
   U307 : BUF_X1 port map( A => n9752, Z => n9755);
   U308 : BUF_X1 port map( A => n9599, Z => n9601);
   U309 : BUF_X1 port map( A => n9598, Z => n9600);
   U310 : BUF_X1 port map( A => n9233, Z => n9599);
   U311 : BUF_X1 port map( A => n9233, Z => n9598);
   U312 : BUF_X1 port map( A => n9233, Z => n9597);
   U313 : BUF_X1 port map( A => n9233, Z => n9596);
   U314 : BUF_X1 port map( A => n9827, Z => n9832);
   U315 : BUF_X1 port map( A => n9826, Z => n9831);
   U316 : BUF_X1 port map( A => n9234, Z => n9830);
   U317 : BUF_X1 port map( A => n9234, Z => n9829);
   U318 : BUF_X1 port map( A => n9234, Z => n9828);
   U319 : BUF_X1 port map( A => n9234, Z => n9827);
   U320 : BUF_X1 port map( A => n9234, Z => n9826);
   U321 : BUF_X1 port map( A => n9234, Z => n9825);
   U322 : BUF_X1 port map( A => n9235, Z => n9715);
   U323 : BUF_X1 port map( A => n9235, Z => n9716);
   U324 : BUF_X1 port map( A => n9235, Z => n9717);
   U325 : BUF_X1 port map( A => n9235, Z => n9718);
   U326 : BUF_X1 port map( A => n9235, Z => n9719);
   U327 : BUF_X1 port map( A => n9235, Z => n9720);
   U328 : BUF_X1 port map( A => n9718, Z => n9721);
   U329 : BUF_X1 port map( A => n9719, Z => n9722);
   U330 : BUF_X1 port map( A => n9629, Z => n9634);
   U331 : BUF_X1 port map( A => n9628, Z => n9633);
   U332 : BUF_X1 port map( A => n9226, Z => n9632);
   U333 : BUF_X1 port map( A => n9226, Z => n9631);
   U334 : BUF_X1 port map( A => n9226, Z => n9630);
   U335 : BUF_X1 port map( A => n9226, Z => n9629);
   U336 : BUF_X1 port map( A => n9226, Z => n9628);
   U337 : BUF_X1 port map( A => n9226, Z => n9627);
   U338 : BUF_X1 port map( A => n9819, Z => n9821);
   U339 : BUF_X1 port map( A => n9818, Z => n9820);
   U340 : BUF_X1 port map( A => n9232, Z => n9819);
   U341 : BUF_X1 port map( A => n9232, Z => n9818);
   U342 : BUF_X1 port map( A => n9232, Z => n9817);
   U343 : BUF_X1 port map( A => n9232, Z => n9816);
   U344 : BUF_X1 port map( A => n9232, Z => n9815);
   U345 : BUF_X1 port map( A => n9232, Z => n9814);
   U346 : BUF_X1 port map( A => n9227, Z => n9693);
   U347 : BUF_X1 port map( A => n9227, Z => n9694);
   U348 : BUF_X1 port map( A => n9227, Z => n9695);
   U349 : BUF_X1 port map( A => n9227, Z => n9696);
   U350 : BUF_X1 port map( A => n9227, Z => n9697);
   U351 : BUF_X1 port map( A => n9227, Z => n9698);
   U352 : BUF_X1 port map( A => n9696, Z => n9699);
   U353 : BUF_X1 port map( A => n9697, Z => n9700);
   U354 : BUF_X1 port map( A => n9805, Z => n9810);
   U355 : BUF_X1 port map( A => n9804, Z => n9809);
   U356 : BUF_X1 port map( A => n9236, Z => n9808);
   U357 : BUF_X1 port map( A => n9236, Z => n9807);
   U358 : BUF_X1 port map( A => n9236, Z => n9806);
   U359 : BUF_X1 port map( A => n9236, Z => n9805);
   U360 : BUF_X1 port map( A => n9236, Z => n9804);
   U361 : BUF_X1 port map( A => n9236, Z => n9803);
   U362 : BUF_X1 port map( A => n9673, Z => n9678);
   U363 : BUF_X1 port map( A => n9672, Z => n9677);
   U364 : BUF_X1 port map( A => n9230, Z => n9676);
   U365 : BUF_X1 port map( A => n9230, Z => n9675);
   U366 : BUF_X1 port map( A => n9230, Z => n9674);
   U367 : BUF_X1 port map( A => n9230, Z => n9673);
   U368 : BUF_X1 port map( A => n9230, Z => n9672);
   U369 : BUF_X1 port map( A => n9230, Z => n9671);
   U370 : BUF_X1 port map( A => n9794, Z => n9799);
   U371 : BUF_X1 port map( A => n9793, Z => n9798);
   U372 : BUF_X1 port map( A => n9237, Z => n9797);
   U373 : BUF_X1 port map( A => n9237, Z => n9796);
   U374 : BUF_X1 port map( A => n9237, Z => n9795);
   U375 : BUF_X1 port map( A => n9237, Z => n9794);
   U376 : BUF_X1 port map( A => n9237, Z => n9793);
   U377 : BUF_X1 port map( A => n9237, Z => n9792);
   U378 : BUF_X1 port map( A => n9884, Z => n9880);
   U379 : BUF_X1 port map( A => n9884, Z => n9882);
   U380 : BUF_X1 port map( A => n9884, Z => n9881);
   U381 : BUF_X1 port map( A => n1516, Z => n9364);
   U382 : BUF_X1 port map( A => n1526, Z => n9340);
   U383 : BUF_X1 port map( A => n1516, Z => n9365);
   U384 : BUF_X1 port map( A => n1526, Z => n9341);
   U385 : BUF_X1 port map( A => n872, Z => n9508);
   U386 : BUF_X1 port map( A => n872, Z => n9509);
   U387 : BUF_X1 port map( A => n877, Z => n9496);
   U388 : BUF_X1 port map( A => n901, Z => n9448);
   U389 : BUF_X1 port map( A => n906, Z => n9436);
   U390 : BUF_X1 port map( A => n882, Z => n9484);
   U391 : BUF_X1 port map( A => n906, Z => n9437);
   U392 : BUF_X1 port map( A => n877, Z => n9497);
   U393 : BUF_X1 port map( A => n867, Z => n9521);
   U394 : BUF_X1 port map( A => n901, Z => n9449);
   U395 : BUF_X1 port map( A => n882, Z => n9485);
   U396 : BUF_X1 port map( A => n1487, Z => n9424);
   U397 : BUF_X1 port map( A => n1492, Z => n9412);
   U398 : BUF_X1 port map( A => n1497, Z => n9400);
   U399 : BUF_X1 port map( A => n1502, Z => n9388);
   U400 : BUF_X1 port map( A => n1511, Z => n9376);
   U401 : BUF_X1 port map( A => n1521, Z => n9352);
   U402 : BUF_X1 port map( A => n1487, Z => n9425);
   U403 : BUF_X1 port map( A => n1492, Z => n9413);
   U404 : BUF_X1 port map( A => n1497, Z => n9401);
   U405 : BUF_X1 port map( A => n1502, Z => n9389);
   U406 : BUF_X1 port map( A => n1511, Z => n9377);
   U407 : BUF_X1 port map( A => n1521, Z => n9353);
   U408 : BUF_X1 port map( A => n893, Z => n9469);
   U409 : BUF_X1 port map( A => n874, Z => n9505);
   U410 : BUF_X1 port map( A => n898, Z => n9457);
   U411 : BUF_X1 port map( A => n884, Z => n9481);
   U412 : BUF_X1 port map( A => n903, Z => n9445);
   U413 : BUF_X1 port map( A => n908, Z => n9433);
   U414 : BUF_X1 port map( A => n879, Z => n9493);
   U415 : BUF_X1 port map( A => n874, Z => n9506);
   U416 : BUF_X1 port map( A => n893, Z => n9470);
   U417 : BUF_X1 port map( A => n898, Z => n9458);
   U418 : BUF_X1 port map( A => n903, Z => n9446);
   U419 : BUF_X1 port map( A => n869, Z => n9518);
   U420 : BUF_X1 port map( A => n884, Z => n9482);
   U421 : BUF_X1 port map( A => n879, Z => n9494);
   U422 : BUF_X1 port map( A => n908, Z => n9434);
   U423 : BUF_X1 port map( A => n1489, Z => n9421);
   U424 : BUF_X1 port map( A => n1494, Z => n9409);
   U425 : BUF_X1 port map( A => n1499, Z => n9397);
   U426 : BUF_X1 port map( A => n1504, Z => n9385);
   U427 : BUF_X1 port map( A => n1513, Z => n9373);
   U428 : BUF_X1 port map( A => n1523, Z => n9349);
   U429 : BUF_X1 port map( A => n1518, Z => n9361);
   U430 : BUF_X1 port map( A => n1528, Z => n9337);
   U431 : BUF_X1 port map( A => n1489, Z => n9422);
   U432 : BUF_X1 port map( A => n1494, Z => n9410);
   U433 : BUF_X1 port map( A => n1499, Z => n9398);
   U434 : BUF_X1 port map( A => n1504, Z => n9386);
   U435 : BUF_X1 port map( A => n1513, Z => n9374);
   U436 : BUF_X1 port map( A => n1523, Z => n9350);
   U437 : BUF_X1 port map( A => n1518, Z => n9362);
   U438 : BUF_X1 port map( A => n1528, Z => n9338);
   U439 : BUF_X1 port map( A => n905, Z => n9439);
   U440 : BUF_X1 port map( A => n905, Z => n9440);
   U441 : BUF_X1 port map( A => n1515, Z => n9367);
   U442 : BUF_X1 port map( A => n1525, Z => n9343);
   U443 : BUF_X1 port map( A => n1515, Z => n9368);
   U444 : BUF_X1 port map( A => n1525, Z => n9344);
   U445 : BUF_X1 port map( A => n871, Z => n9511);
   U446 : BUF_X1 port map( A => n871, Z => n9512);
   U447 : BUF_X1 port map( A => n1491, Z => n9415);
   U448 : BUF_X1 port map( A => n1491, Z => n9416);
   U449 : BUF_X1 port map( A => n900, Z => n9451);
   U450 : BUF_X1 port map( A => n876, Z => n9499);
   U451 : BUF_X1 port map( A => n881, Z => n9487);
   U452 : BUF_X1 port map( A => n866, Z => n9524);
   U453 : BUF_X1 port map( A => n900, Z => n9452);
   U454 : BUF_X1 port map( A => n876, Z => n9500);
   U455 : BUF_X1 port map( A => n881, Z => n9488);
   U456 : BUF_X1 port map( A => n1486, Z => n9427);
   U457 : BUF_X1 port map( A => n1496, Z => n9403);
   U458 : BUF_X1 port map( A => n1501, Z => n9391);
   U459 : BUF_X1 port map( A => n1510, Z => n9379);
   U460 : BUF_X1 port map( A => n1520, Z => n9355);
   U461 : BUF_X1 port map( A => n1486, Z => n9428);
   U462 : BUF_X1 port map( A => n1496, Z => n9404);
   U463 : BUF_X1 port map( A => n1501, Z => n9392);
   U464 : BUF_X1 port map( A => n1510, Z => n9380);
   U465 : BUF_X1 port map( A => n1520, Z => n9356);
   U466 : BUF_X1 port map( A => n867, Z => n9520);
   U467 : BUF_X1 port map( A => n869, Z => n9517);
   U468 : BUF_X1 port map( A => n866, Z => n9523);
   U469 : BUF_X1 port map( A => n885, Z => n9478);
   U470 : BUF_X1 port map( A => n894, Z => n9466);
   U471 : BUF_X1 port map( A => n870, Z => n9514);
   U472 : BUF_X1 port map( A => n899, Z => n9454);
   U473 : BUF_X1 port map( A => n880, Z => n9490);
   U474 : BUF_X1 port map( A => n875, Z => n9502);
   U475 : BUF_X1 port map( A => n904, Z => n9442);
   U476 : BUF_X1 port map( A => n875, Z => n9503);
   U477 : BUF_X1 port map( A => n870, Z => n9515);
   U478 : BUF_X1 port map( A => n894, Z => n9467);
   U479 : BUF_X1 port map( A => n899, Z => n9455);
   U480 : BUF_X1 port map( A => n885, Z => n9479);
   U481 : BUF_X1 port map( A => n880, Z => n9491);
   U482 : BUF_X1 port map( A => n904, Z => n9443);
   U483 : BUF_X1 port map( A => n909, Z => n9430);
   U484 : BUF_X1 port map( A => n909, Z => n9431);
   U485 : BUF_X1 port map( A => n1490, Z => n9419);
   U486 : BUF_X1 port map( A => n1495, Z => n9407);
   U487 : BUF_X1 port map( A => n1500, Z => n9395);
   U488 : BUF_X1 port map( A => n1505, Z => n9383);
   U489 : BUF_X1 port map( A => n1514, Z => n9371);
   U490 : BUF_X1 port map( A => n1524, Z => n9347);
   U491 : BUF_X1 port map( A => n1519, Z => n9359);
   U492 : BUF_X1 port map( A => n1529, Z => n9335);
   U493 : BUF_X1 port map( A => n1490, Z => n9418);
   U494 : BUF_X1 port map( A => n1495, Z => n9406);
   U495 : BUF_X1 port map( A => n1500, Z => n9394);
   U496 : BUF_X1 port map( A => n1505, Z => n9382);
   U497 : BUF_X1 port map( A => n1514, Z => n9370);
   U498 : BUF_X1 port map( A => n1524, Z => n9346);
   U499 : BUF_X1 port map( A => n1519, Z => n9358);
   U500 : BUF_X1 port map( A => n1529, Z => n9334);
   U501 : BUF_X1 port map( A => n891, Z => n9472);
   U502 : BUF_X1 port map( A => n896, Z => n9460);
   U503 : BUF_X1 port map( A => n896, Z => n9461);
   U504 : BUF_X1 port map( A => n891, Z => n9473);
   U505 : BUF_X1 port map( A => n1516, Z => n9366);
   U506 : BUF_X1 port map( A => n1526, Z => n9342);
   U507 : BUF_X1 port map( A => n1492, Z => n9414);
   U508 : BUF_X1 port map( A => n882, Z => n9486);
   U509 : BUF_X1 port map( A => n867, Z => n9522);
   U510 : BUF_X1 port map( A => n877, Z => n9498);
   U511 : BUF_X1 port map( A => n896, Z => n9462);
   U512 : BUF_X1 port map( A => n891, Z => n9474);
   U513 : BUF_X1 port map( A => n901, Z => n9450);
   U514 : BUF_X1 port map( A => n872, Z => n9510);
   U515 : BUF_X1 port map( A => n906, Z => n9438);
   U516 : BUF_X1 port map( A => n1487, Z => n9426);
   U517 : BUF_X1 port map( A => n1497, Z => n9402);
   U518 : BUF_X1 port map( A => n1502, Z => n9390);
   U519 : BUF_X1 port map( A => n1511, Z => n9378);
   U520 : BUF_X1 port map( A => n1521, Z => n9354);
   U521 : BUF_X1 port map( A => n890, Z => n9475);
   U522 : BUF_X1 port map( A => n895, Z => n9463);
   U523 : BUF_X1 port map( A => n890, Z => n9476);
   U524 : BUF_X1 port map( A => n895, Z => n9464);
   U525 : BUF_X1 port map( A => n898, Z => n9459);
   U526 : BUF_X1 port map( A => n869, Z => n9519);
   U527 : BUF_X1 port map( A => n893, Z => n9471);
   U528 : BUF_X1 port map( A => n884, Z => n9483);
   U529 : BUF_X1 port map( A => n903, Z => n9447);
   U530 : BUF_X1 port map( A => n874, Z => n9507);
   U531 : BUF_X1 port map( A => n879, Z => n9495);
   U532 : BUF_X1 port map( A => n908, Z => n9435);
   U533 : BUF_X1 port map( A => n1489, Z => n9423);
   U534 : BUF_X1 port map( A => n1494, Z => n9411);
   U535 : BUF_X1 port map( A => n1499, Z => n9399);
   U536 : BUF_X1 port map( A => n1504, Z => n9387);
   U537 : BUF_X1 port map( A => n1513, Z => n9375);
   U538 : BUF_X1 port map( A => n1523, Z => n9351);
   U539 : BUF_X1 port map( A => n1518, Z => n9363);
   U540 : BUF_X1 port map( A => n1528, Z => n9339);
   U541 : BUF_X1 port map( A => n905, Z => n9441);
   U542 : BUF_X1 port map( A => n1515, Z => n9369);
   U543 : BUF_X1 port map( A => n1525, Z => n9345);
   U544 : BUF_X1 port map( A => n1491, Z => n9417);
   U545 : BUF_X1 port map( A => n881, Z => n9489);
   U546 : BUF_X1 port map( A => n890, Z => n9477);
   U547 : BUF_X1 port map( A => n866, Z => n9525);
   U548 : BUF_X1 port map( A => n895, Z => n9465);
   U549 : BUF_X1 port map( A => n871, Z => n9513);
   U550 : BUF_X1 port map( A => n900, Z => n9453);
   U551 : BUF_X1 port map( A => n876, Z => n9501);
   U552 : BUF_X1 port map( A => n1486, Z => n9429);
   U553 : BUF_X1 port map( A => n1496, Z => n9405);
   U554 : BUF_X1 port map( A => n1501, Z => n9393);
   U555 : BUF_X1 port map( A => n1510, Z => n9381);
   U556 : BUF_X1 port map( A => n1520, Z => n9357);
   U557 : BUF_X1 port map( A => n875, Z => n9504);
   U558 : BUF_X1 port map( A => n885, Z => n9480);
   U559 : BUF_X1 port map( A => n899, Z => n9456);
   U560 : BUF_X1 port map( A => n909, Z => n9432);
   U561 : BUF_X1 port map( A => n894, Z => n9468);
   U562 : BUF_X1 port map( A => n880, Z => n9492);
   U563 : BUF_X1 port map( A => n904, Z => n9444);
   U564 : BUF_X1 port map( A => n1514, Z => n9372);
   U565 : BUF_X1 port map( A => n1524, Z => n9348);
   U566 : BUF_X1 port map( A => n1519, Z => n9360);
   U567 : BUF_X1 port map( A => n1529, Z => n9336);
   U568 : BUF_X1 port map( A => n1490, Z => n9420);
   U569 : BUF_X1 port map( A => n1495, Z => n9408);
   U570 : BUF_X1 port map( A => n1500, Z => n9396);
   U571 : BUF_X1 port map( A => n1505, Z => n9384);
   U572 : BUF_X1 port map( A => n870, Z => n9516);
   U573 : BUF_X1 port map( A => n815, Z => n9874);
   U574 : BUF_X1 port map( A => n815, Z => n9873);
   U575 : BUF_X1 port map( A => n815, Z => n9872);
   U576 : BUF_X1 port map( A => n815, Z => n9871);
   U577 : BUF_X1 port map( A => n815, Z => n9870);
   U578 : BUF_X1 port map( A => n815, Z => n9869);
   U579 : BUF_X1 port map( A => n815, Z => n9875);
   U580 : INV_X1 port map( A => n9876, ZN => n9884);
   U581 : NOR3_X1 port map( A1 => n9920, A2 => n9919, A3 => n9921, ZN => n824);
   U582 : AND3_X1 port map( A1 => n9918, A2 => n9917, A3 => n849, ZN => n830);
   U583 : BUF_X1 port map( A => n9916, Z => n9331);
   U584 : BUF_X1 port map( A => n9915, Z => n9328);
   U585 : BUF_X1 port map( A => n9914, Z => n9325);
   U586 : BUF_X1 port map( A => n9913, Z => n9322);
   U587 : BUF_X1 port map( A => n9912, Z => n9319);
   U588 : BUF_X1 port map( A => n9911, Z => n9316);
   U589 : BUF_X1 port map( A => n9910, Z => n9313);
   U590 : BUF_X1 port map( A => n9909, Z => n9310);
   U591 : BUF_X1 port map( A => n9908, Z => n9307);
   U592 : BUF_X1 port map( A => n9907, Z => n9304);
   U593 : BUF_X1 port map( A => n9906, Z => n9301);
   U594 : BUF_X1 port map( A => n9905, Z => n9298);
   U595 : BUF_X1 port map( A => n9904, Z => n9295);
   U596 : BUF_X1 port map( A => n9903, Z => n9292);
   U597 : BUF_X1 port map( A => n9902, Z => n9289);
   U598 : BUF_X1 port map( A => n9901, Z => n9286);
   U599 : BUF_X1 port map( A => n9900, Z => n9283);
   U600 : BUF_X1 port map( A => n9899, Z => n9280);
   U601 : BUF_X1 port map( A => n9898, Z => n9277);
   U602 : BUF_X1 port map( A => n9897, Z => n9274);
   U603 : BUF_X1 port map( A => n9896, Z => n9271);
   U604 : BUF_X1 port map( A => n9895, Z => n9268);
   U605 : BUF_X1 port map( A => n9894, Z => n9265);
   U606 : BUF_X1 port map( A => n9893, Z => n9262);
   U607 : BUF_X1 port map( A => n9892, Z => n9259);
   U608 : BUF_X1 port map( A => n9891, Z => n9256);
   U609 : BUF_X1 port map( A => n9890, Z => n9253);
   U610 : BUF_X1 port map( A => n9889, Z => n9250);
   U611 : BUF_X1 port map( A => n9888, Z => n9247);
   U612 : BUF_X1 port map( A => n9887, Z => n9244);
   U613 : BUF_X1 port map( A => n9886, Z => n9241);
   U614 : BUF_X1 port map( A => n9885, Z => n9238);
   U615 : BUF_X1 port map( A => n9916, Z => n9332);
   U616 : BUF_X1 port map( A => n9915, Z => n9329);
   U617 : BUF_X1 port map( A => n9914, Z => n9326);
   U618 : BUF_X1 port map( A => n9913, Z => n9323);
   U619 : BUF_X1 port map( A => n9912, Z => n9320);
   U620 : BUF_X1 port map( A => n9911, Z => n9317);
   U621 : BUF_X1 port map( A => n9910, Z => n9314);
   U622 : BUF_X1 port map( A => n9909, Z => n9311);
   U623 : BUF_X1 port map( A => n9908, Z => n9308);
   U624 : BUF_X1 port map( A => n9907, Z => n9305);
   U625 : BUF_X1 port map( A => n9906, Z => n9302);
   U626 : BUF_X1 port map( A => n9905, Z => n9299);
   U627 : BUF_X1 port map( A => n9904, Z => n9296);
   U628 : BUF_X1 port map( A => n9903, Z => n9293);
   U629 : BUF_X1 port map( A => n9902, Z => n9290);
   U630 : BUF_X1 port map( A => n9901, Z => n9287);
   U631 : BUF_X1 port map( A => n9900, Z => n9284);
   U632 : BUF_X1 port map( A => n9899, Z => n9281);
   U633 : BUF_X1 port map( A => n9898, Z => n9278);
   U634 : BUF_X1 port map( A => n9897, Z => n9275);
   U635 : BUF_X1 port map( A => n9896, Z => n9272);
   U636 : BUF_X1 port map( A => n9895, Z => n9269);
   U637 : BUF_X1 port map( A => n9894, Z => n9266);
   U638 : BUF_X1 port map( A => n9893, Z => n9263);
   U639 : BUF_X1 port map( A => n9892, Z => n9260);
   U640 : BUF_X1 port map( A => n9891, Z => n9257);
   U641 : BUF_X1 port map( A => n9890, Z => n9254);
   U642 : BUF_X1 port map( A => n9889, Z => n9251);
   U643 : BUF_X1 port map( A => n9888, Z => n9248);
   U644 : BUF_X1 port map( A => n9887, Z => n9245);
   U645 : BUF_X1 port map( A => n9886, Z => n9242);
   U646 : BUF_X1 port map( A => n9885, Z => n9239);
   U647 : NAND2_X1 port map( A1 => n1459, A2 => n1458, ZN => n866);
   U648 : NAND2_X1 port map( A1 => n1457, A2 => n1470, ZN => n896);
   U649 : AOI22_X1 port map( A1 => n9483, A2 => n10194, B1 => n9478, B2 => 
                           n10554, ZN => n883);
   U650 : AOI22_X1 port map( A1 => n9483, A2 => n10200, B1 => n9478, B2 => 
                           n10560, ZN => n1009);
   U651 : AOI22_X1 port map( A1 => n9483, A2 => n10197, B1 => n9478, B2 => 
                           n10557, ZN => n955);
   U652 : AOI22_X1 port map( A1 => n9483, A2 => n10201, B1 => n9478, B2 => 
                           n10561, ZN => n1027);
   U653 : AOI22_X1 port map( A1 => n9483, A2 => n10196, B1 => n9478, B2 => 
                           n10556, ZN => n937);
   U654 : AOI22_X1 port map( A1 => n9483, A2 => n10199, B1 => n9478, B2 => 
                           n10559, ZN => n991);
   U655 : AOI22_X1 port map( A1 => n9483, A2 => n10195, B1 => n9478, B2 => 
                           n10555, ZN => n919);
   U656 : AOI22_X1 port map( A1 => n9483, A2 => n10198, B1 => n9478, B2 => 
                           n10558, ZN => n973);
   U657 : NAND2_X1 port map( A1 => n2084, A2 => n2088, ZN => n1501);
   U658 : NAND2_X1 port map( A1 => n2083, A2 => n2088, ZN => n1502);
   U659 : NAND2_X1 port map( A1 => n1477, A2 => n1459, ZN => n905);
   U660 : NAND2_X1 port map( A1 => n1461, A2 => n1460, ZN => n872);
   U661 : NAND2_X1 port map( A1 => n1461, A2 => n1458, ZN => n867);
   U662 : NAND2_X1 port map( A1 => n816, A2 => n817, ZN => n815);
   U663 : BUF_X1 port map( A => n9916, Z => n9333);
   U664 : BUF_X1 port map( A => n9915, Z => n9330);
   U665 : BUF_X1 port map( A => n9914, Z => n9327);
   U666 : BUF_X1 port map( A => n9913, Z => n9324);
   U667 : BUF_X1 port map( A => n9912, Z => n9321);
   U668 : BUF_X1 port map( A => n9911, Z => n9318);
   U669 : BUF_X1 port map( A => n9910, Z => n9315);
   U670 : BUF_X1 port map( A => n9909, Z => n9312);
   U671 : BUF_X1 port map( A => n9908, Z => n9309);
   U672 : BUF_X1 port map( A => n9907, Z => n9306);
   U673 : BUF_X1 port map( A => n9906, Z => n9303);
   U674 : BUF_X1 port map( A => n9905, Z => n9300);
   U675 : BUF_X1 port map( A => n9904, Z => n9297);
   U676 : BUF_X1 port map( A => n9903, Z => n9294);
   U677 : BUF_X1 port map( A => n9902, Z => n9291);
   U678 : BUF_X1 port map( A => n9901, Z => n9288);
   U679 : BUF_X1 port map( A => n9900, Z => n9285);
   U680 : BUF_X1 port map( A => n9899, Z => n9282);
   U681 : BUF_X1 port map( A => n9898, Z => n9279);
   U682 : BUF_X1 port map( A => n9897, Z => n9276);
   U683 : BUF_X1 port map( A => n9896, Z => n9273);
   U684 : BUF_X1 port map( A => n9895, Z => n9270);
   U685 : BUF_X1 port map( A => n9894, Z => n9267);
   U686 : BUF_X1 port map( A => n9893, Z => n9264);
   U687 : BUF_X1 port map( A => n9892, Z => n9261);
   U688 : BUF_X1 port map( A => n9891, Z => n9258);
   U689 : BUF_X1 port map( A => n9890, Z => n9255);
   U690 : BUF_X1 port map( A => n9889, Z => n9252);
   U691 : BUF_X1 port map( A => n9888, Z => n9249);
   U692 : BUF_X1 port map( A => n9887, Z => n9246);
   U693 : BUF_X1 port map( A => n9886, Z => n9243);
   U694 : BUF_X1 port map( A => n9885, Z => n9240);
   U695 : NAND2_X1 port map( A1 => n2095, A2 => n2084, ZN => n1515);
   U696 : NAND2_X1 port map( A1 => n2095, A2 => n2083, ZN => n1516);
   U697 : NAND2_X1 port map( A1 => n2098, A2 => n2084, ZN => n1525);
   U698 : NAND2_X1 port map( A1 => n2098, A2 => n2083, ZN => n1526);
   U699 : NAND2_X1 port map( A1 => n1477, A2 => n1461, ZN => n906);
   U700 : NAND2_X1 port map( A1 => n1464, A2 => n1460, ZN => n881);
   U701 : NAND2_X1 port map( A1 => n2077, A2 => n2085, ZN => n1492);
   U702 : NAND2_X1 port map( A1 => n2077, A2 => n2086, ZN => n1491);
   U703 : NAND2_X1 port map( A1 => n1458, A2 => n1464, ZN => n871);
   U704 : NAND2_X1 port map( A1 => n1470, A2 => n1464, ZN => n891);
   U705 : NAND2_X1 port map( A1 => n1477, A2 => n1464, ZN => n895);
   U706 : NAND2_X1 port map( A1 => n1468, A2 => n1470, ZN => n890);
   U707 : AND2_X1 port map( A1 => n1459, A2 => n1470, ZN => n898);
   U708 : AND2_X1 port map( A1 => n1459, A2 => n1460, ZN => n869);
   U709 : NAND2_X1 port map( A1 => n1458, A2 => n1468, ZN => n877);
   U710 : NAND2_X1 port map( A1 => n1477, A2 => n1468, ZN => n901);
   U711 : NAND2_X1 port map( A1 => n1458, A2 => n1467, ZN => n876);
   U712 : NAND2_X1 port map( A1 => n2079, A2 => n2088, ZN => n1496);
   U713 : NAND2_X1 port map( A1 => n2078, A2 => n2088, ZN => n1497);
   U714 : AND2_X1 port map( A1 => n1457, A2 => n1460, ZN => n875);
   U715 : AND2_X1 port map( A1 => n1457, A2 => n1458, ZN => n870);
   U716 : NAND2_X1 port map( A1 => n1466, A2 => n1460, ZN => n882);
   U717 : NAND2_X1 port map( A1 => n2095, A2 => n2079, ZN => n1510);
   U718 : NAND2_X1 port map( A1 => n2095, A2 => n2078, ZN => n1511);
   U719 : NAND2_X1 port map( A1 => n2098, A2 => n2079, ZN => n1520);
   U720 : NAND2_X1 port map( A1 => n2098, A2 => n2078, ZN => n1521);
   U721 : NAND2_X1 port map( A1 => n1477, A2 => n1467, ZN => n900);
   U722 : NAND2_X1 port map( A1 => n2077, A2 => n2081, ZN => n1486);
   U723 : NAND2_X1 port map( A1 => n2077, A2 => n2080, ZN => n1487);
   U724 : AND2_X1 port map( A1 => n1477, A2 => n1457, ZN => n909);
   U725 : AND2_X1 port map( A1 => n1461, A2 => n1470, ZN => n899);
   U726 : AND2_X1 port map( A1 => n2085, A2 => n2088, ZN => n1505);
   U727 : AND2_X1 port map( A1 => n2086, A2 => n2088, ZN => n1504);
   U728 : AND2_X1 port map( A1 => n2077, A2 => n2083, ZN => n1495);
   U729 : AND2_X1 port map( A1 => n2077, A2 => n2084, ZN => n1494);
   U730 : AND2_X1 port map( A1 => n1463, A2 => n1470, ZN => n893);
   U731 : AND2_X1 port map( A1 => n1463, A2 => n1460, ZN => n874);
   U732 : AND2_X1 port map( A1 => n1463, A2 => n1458, ZN => n908);
   U733 : AND2_X1 port map( A1 => n2095, A2 => n2085, ZN => n1519);
   U734 : AND2_X1 port map( A1 => n2095, A2 => n2086, ZN => n1518);
   U735 : AND2_X1 port map( A1 => n2098, A2 => n2085, ZN => n1529);
   U736 : AND2_X1 port map( A1 => n2098, A2 => n2086, ZN => n1528);
   U737 : AND2_X1 port map( A1 => n1477, A2 => n1463, ZN => n903);
   U738 : AND2_X1 port map( A1 => n1468, A2 => n1460, ZN => n885);
   U739 : AND2_X1 port map( A1 => n1458, A2 => n1466, ZN => n880);
   U740 : AND2_X1 port map( A1 => n1477, A2 => n1466, ZN => n904);
   U741 : AND2_X1 port map( A1 => n2077, A2 => n2079, ZN => n1489);
   U742 : AND2_X1 port map( A1 => n2077, A2 => n2078, ZN => n1490);
   U743 : AND2_X1 port map( A1 => n2095, A2 => n2081, ZN => n1513);
   U744 : AND2_X1 port map( A1 => n2095, A2 => n2080, ZN => n1514);
   U745 : AND2_X1 port map( A1 => n2098, A2 => n2081, ZN => n1523);
   U746 : AND2_X1 port map( A1 => n2098, A2 => n2080, ZN => n1524);
   U747 : AND2_X1 port map( A1 => n1470, A2 => n1466, ZN => n884);
   U748 : AND2_X1 port map( A1 => n2081, A2 => n2088, ZN => n1499);
   U749 : AND2_X1 port map( A1 => n2080, A2 => n2088, ZN => n1500);
   U750 : AND2_X1 port map( A1 => n1467, A2 => n1460, ZN => n879);
   U751 : AND2_X1 port map( A1 => n1467, A2 => n1470, ZN => n894);
   U752 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(1), A3 => n9919, ZN 
                           => n817);
   U753 : NOR3_X1 port map( A1 => ADD_WR(0), A2 => ADD_WR(2), A3 => n9920, ZN 
                           => n822);
   U754 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => ADD_WR(0), 
                           ZN => n819);
   U755 : NOR3_X1 port map( A1 => n9919, A2 => ADD_WR(1), A3 => n9921, ZN => 
                           n827);
   U756 : NOR3_X1 port map( A1 => n9919, A2 => ADD_WR(0), A3 => n9920, ZN => 
                           n847);
   U757 : NOR3_X1 port map( A1 => n9920, A2 => ADD_WR(2), A3 => n9921, ZN => 
                           n845);
   U758 : NOR3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(2), A3 => n9921, ZN 
                           => n842);
   U759 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(2), A3 => n10663, 
                           ZN => n2084);
   U760 : NOR3_X1 port map( A1 => n10664, A2 => ADD_RD2(2), A3 => n10663, ZN =>
                           n2083);
   U761 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(2), A3 => n10659, 
                           ZN => n1461);
   U762 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n10664, 
                           ZN => n2085);
   U763 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => 
                           ADD_RD2(0), ZN => n2086);
   U764 : NOR3_X1 port map( A1 => n10660, A2 => ADD_RD1(2), A3 => n10659, ZN =>
                           n1463);
   U765 : NOR4_X1 port map( A1 => n1928, A2 => n1929, A3 => n1930, A4 => n1931,
                           ZN => n1927);
   U766 : OAI221_X1 port map( B1 => n8574, B2 => n9391, C1 => n8550, C2 => 
                           n9388, A => n1935, ZN => n1928);
   U767 : OAI221_X1 port map( B1 => n8486, B2 => n9403, C1 => n8247, C2 => 
                           n9400, A => n1934, ZN => n1929);
   U768 : OAI221_X1 port map( B1 => n8447, B2 => n9415, C1 => n8415, C2 => 
                           n9412, A => n1933, ZN => n1930);
   U769 : NOR4_X1 port map( A1 => n1910, A2 => n1911, A3 => n1912, A4 => n1913,
                           ZN => n1909);
   U770 : OAI221_X1 port map( B1 => n8575, B2 => n9391, C1 => n8551, C2 => 
                           n9388, A => n1917, ZN => n1910);
   U771 : OAI221_X1 port map( B1 => n8487, B2 => n9403, C1 => n8248, C2 => 
                           n9400, A => n1916, ZN => n1911);
   U772 : OAI221_X1 port map( B1 => n8448, B2 => n9415, C1 => n8416, C2 => 
                           n9412, A => n1915, ZN => n1912);
   U773 : NOR4_X1 port map( A1 => n1892, A2 => n1893, A3 => n1894, A4 => n1895,
                           ZN => n1891);
   U774 : OAI221_X1 port map( B1 => n8576, B2 => n9391, C1 => n8552, C2 => 
                           n9388, A => n1899, ZN => n1892);
   U775 : OAI221_X1 port map( B1 => n8488, B2 => n9403, C1 => n8249, C2 => 
                           n9400, A => n1898, ZN => n1893);
   U776 : OAI221_X1 port map( B1 => n8449, B2 => n9415, C1 => n8417, C2 => 
                           n9412, A => n1897, ZN => n1894);
   U777 : NOR4_X1 port map( A1 => n1874, A2 => n1875, A3 => n1876, A4 => n1877,
                           ZN => n1873);
   U778 : OAI221_X1 port map( B1 => n8577, B2 => n9391, C1 => n8553, C2 => 
                           n9388, A => n1881, ZN => n1874);
   U779 : OAI221_X1 port map( B1 => n8489, B2 => n9403, C1 => n8250, C2 => 
                           n9400, A => n1880, ZN => n1875);
   U780 : OAI221_X1 port map( B1 => n8450, B2 => n9415, C1 => n8418, C2 => 
                           n9412, A => n1879, ZN => n1876);
   U781 : NOR4_X1 port map( A1 => n1856, A2 => n1857, A3 => n1858, A4 => n1859,
                           ZN => n1855);
   U782 : OAI221_X1 port map( B1 => n8578, B2 => n9392, C1 => n8554, C2 => 
                           n9389, A => n1863, ZN => n1856);
   U783 : OAI221_X1 port map( B1 => n8490, B2 => n9404, C1 => n8251, C2 => 
                           n9401, A => n1862, ZN => n1857);
   U784 : OAI221_X1 port map( B1 => n8451, B2 => n9416, C1 => n8419, C2 => 
                           n9413, A => n1861, ZN => n1858);
   U785 : NOR4_X1 port map( A1 => n1838, A2 => n1839, A3 => n1840, A4 => n1841,
                           ZN => n1837);
   U786 : OAI221_X1 port map( B1 => n8579, B2 => n9392, C1 => n8555, C2 => 
                           n9389, A => n1845, ZN => n1838);
   U787 : OAI221_X1 port map( B1 => n8491, B2 => n9404, C1 => n8252, C2 => 
                           n9401, A => n1844, ZN => n1839);
   U788 : OAI221_X1 port map( B1 => n8452, B2 => n9416, C1 => n8420, C2 => 
                           n9413, A => n1843, ZN => n1840);
   U789 : NOR4_X1 port map( A1 => n1820, A2 => n1821, A3 => n1822, A4 => n1823,
                           ZN => n1819);
   U790 : OAI221_X1 port map( B1 => n8580, B2 => n9392, C1 => n8556, C2 => 
                           n9389, A => n1827, ZN => n1820);
   U791 : OAI221_X1 port map( B1 => n8492, B2 => n9404, C1 => n8253, C2 => 
                           n9401, A => n1826, ZN => n1821);
   U792 : OAI221_X1 port map( B1 => n8453, B2 => n9416, C1 => n8421, C2 => 
                           n9413, A => n1825, ZN => n1822);
   U793 : NOR4_X1 port map( A1 => n1802, A2 => n1803, A3 => n1804, A4 => n1805,
                           ZN => n1801);
   U794 : OAI221_X1 port map( B1 => n8581, B2 => n9392, C1 => n8557, C2 => 
                           n9389, A => n1809, ZN => n1802);
   U795 : OAI221_X1 port map( B1 => n8493, B2 => n9404, C1 => n8254, C2 => 
                           n9401, A => n1808, ZN => n1803);
   U796 : OAI221_X1 port map( B1 => n8454, B2 => n9416, C1 => n8422, C2 => 
                           n9413, A => n1807, ZN => n1804);
   U797 : NOR4_X1 port map( A1 => n1784, A2 => n1785, A3 => n1786, A4 => n1787,
                           ZN => n1783);
   U798 : OAI221_X1 port map( B1 => n8582, B2 => n9392, C1 => n8558, C2 => 
                           n9389, A => n1791, ZN => n1784);
   U799 : OAI221_X1 port map( B1 => n8494, B2 => n9404, C1 => n8255, C2 => 
                           n9401, A => n1790, ZN => n1785);
   U800 : OAI221_X1 port map( B1 => n8455, B2 => n9416, C1 => n8423, C2 => 
                           n9413, A => n1789, ZN => n1786);
   U801 : NOR4_X1 port map( A1 => n1766, A2 => n1767, A3 => n1768, A4 => n1769,
                           ZN => n1765);
   U802 : OAI221_X1 port map( B1 => n8583, B2 => n9392, C1 => n8559, C2 => 
                           n9389, A => n1773, ZN => n1766);
   U803 : OAI221_X1 port map( B1 => n8495, B2 => n9404, C1 => n8256, C2 => 
                           n9401, A => n1772, ZN => n1767);
   U804 : OAI221_X1 port map( B1 => n8456, B2 => n9416, C1 => n8424, C2 => 
                           n9413, A => n1771, ZN => n1768);
   U805 : NOR4_X1 port map( A1 => n1748, A2 => n1749, A3 => n1750, A4 => n1751,
                           ZN => n1747);
   U806 : OAI221_X1 port map( B1 => n8584, B2 => n9392, C1 => n8560, C2 => 
                           n9389, A => n1755, ZN => n1748);
   U807 : OAI221_X1 port map( B1 => n8496, B2 => n9404, C1 => n8257, C2 => 
                           n9401, A => n1754, ZN => n1749);
   U808 : OAI221_X1 port map( B1 => n8457, B2 => n9416, C1 => n8425, C2 => 
                           n9413, A => n1753, ZN => n1750);
   U809 : NOR4_X1 port map( A1 => n1730, A2 => n1731, A3 => n1732, A4 => n1733,
                           ZN => n1729);
   U810 : OAI221_X1 port map( B1 => n8585, B2 => n9392, C1 => n8561, C2 => 
                           n9389, A => n1737, ZN => n1730);
   U811 : OAI221_X1 port map( B1 => n8497, B2 => n9404, C1 => n8258, C2 => 
                           n9401, A => n1736, ZN => n1731);
   U812 : OAI221_X1 port map( B1 => n8458, B2 => n9416, C1 => n8426, C2 => 
                           n9413, A => n1735, ZN => n1732);
   U813 : NOR4_X1 port map( A1 => n1712, A2 => n1713, A3 => n1714, A4 => n1715,
                           ZN => n1711);
   U814 : OAI221_X1 port map( B1 => n8586, B2 => n9392, C1 => n8562, C2 => 
                           n9389, A => n1719, ZN => n1712);
   U815 : OAI221_X1 port map( B1 => n8498, B2 => n9404, C1 => n8259, C2 => 
                           n9401, A => n1718, ZN => n1713);
   U816 : OAI221_X1 port map( B1 => n8459, B2 => n9416, C1 => n8427, C2 => 
                           n9413, A => n1717, ZN => n1714);
   U817 : NOR4_X1 port map( A1 => n1694, A2 => n1695, A3 => n1696, A4 => n1697,
                           ZN => n1693);
   U818 : OAI221_X1 port map( B1 => n8587, B2 => n9392, C1 => n8563, C2 => 
                           n9389, A => n1701, ZN => n1694);
   U819 : OAI221_X1 port map( B1 => n8499, B2 => n9404, C1 => n8260, C2 => 
                           n9401, A => n1700, ZN => n1695);
   U820 : OAI221_X1 port map( B1 => n8460, B2 => n9416, C1 => n8428, C2 => 
                           n9413, A => n1699, ZN => n1696);
   U821 : NOR4_X1 port map( A1 => n1676, A2 => n1677, A3 => n1678, A4 => n1679,
                           ZN => n1675);
   U822 : OAI221_X1 port map( B1 => n8588, B2 => n9392, C1 => n8564, C2 => 
                           n9389, A => n1683, ZN => n1676);
   U823 : OAI221_X1 port map( B1 => n8500, B2 => n9404, C1 => n8261, C2 => 
                           n9401, A => n1682, ZN => n1677);
   U824 : OAI221_X1 port map( B1 => n8461, B2 => n9416, C1 => n8429, C2 => 
                           n9413, A => n1681, ZN => n1678);
   U825 : NOR4_X1 port map( A1 => n1658, A2 => n1659, A3 => n1660, A4 => n1661,
                           ZN => n1657);
   U826 : OAI221_X1 port map( B1 => n8589, B2 => n9392, C1 => n8565, C2 => 
                           n9389, A => n1665, ZN => n1658);
   U827 : OAI221_X1 port map( B1 => n8501, B2 => n9404, C1 => n8262, C2 => 
                           n9401, A => n1664, ZN => n1659);
   U828 : OAI221_X1 port map( B1 => n8462, B2 => n9416, C1 => n8430, C2 => 
                           n9413, A => n1663, ZN => n1660);
   U829 : NOR4_X1 port map( A1 => n1640, A2 => n1641, A3 => n1642, A4 => n1643,
                           ZN => n1639);
   U830 : OAI221_X1 port map( B1 => n8590, B2 => n9393, C1 => n8319, C2 => 
                           n9390, A => n1647, ZN => n1640);
   U831 : OAI221_X1 port map( B1 => n8502, B2 => n9405, C1 => n8327, C2 => 
                           n9402, A => n1646, ZN => n1641);
   U832 : OAI221_X1 port map( B1 => n8463, B2 => n9417, C1 => n8431, C2 => 
                           n9414, A => n1645, ZN => n1642);
   U833 : NOR4_X1 port map( A1 => n1622, A2 => n1623, A3 => n1624, A4 => n1625,
                           ZN => n1621);
   U834 : OAI221_X1 port map( B1 => n8591, B2 => n9393, C1 => n8320, C2 => 
                           n9390, A => n1629, ZN => n1622);
   U835 : OAI221_X1 port map( B1 => n8503, B2 => n9405, C1 => n8328, C2 => 
                           n9402, A => n1628, ZN => n1623);
   U836 : OAI221_X1 port map( B1 => n8464, B2 => n9417, C1 => n8432, C2 => 
                           n9414, A => n1627, ZN => n1624);
   U837 : NOR4_X1 port map( A1 => n1604, A2 => n1605, A3 => n1606, A4 => n1607,
                           ZN => n1603);
   U838 : OAI221_X1 port map( B1 => n8592, B2 => n9393, C1 => n8321, C2 => 
                           n9390, A => n1611, ZN => n1604);
   U839 : OAI221_X1 port map( B1 => n8504, B2 => n9405, C1 => n8329, C2 => 
                           n9402, A => n1610, ZN => n1605);
   U840 : OAI221_X1 port map( B1 => n8465, B2 => n9417, C1 => n8433, C2 => 
                           n9414, A => n1609, ZN => n1606);
   U841 : NOR4_X1 port map( A1 => n1586, A2 => n1587, A3 => n1588, A4 => n1589,
                           ZN => n1585);
   U842 : OAI221_X1 port map( B1 => n8593, B2 => n9393, C1 => n8322, C2 => 
                           n9390, A => n1593, ZN => n1586);
   U843 : OAI221_X1 port map( B1 => n8505, B2 => n9405, C1 => n8330, C2 => 
                           n9402, A => n1592, ZN => n1587);
   U844 : OAI221_X1 port map( B1 => n8466, B2 => n9417, C1 => n8434, C2 => 
                           n9414, A => n1591, ZN => n1588);
   U845 : NOR4_X1 port map( A1 => n1568, A2 => n1569, A3 => n1570, A4 => n1571,
                           ZN => n1567);
   U846 : OAI221_X1 port map( B1 => n8594, B2 => n9393, C1 => n8323, C2 => 
                           n9390, A => n1575, ZN => n1568);
   U847 : OAI221_X1 port map( B1 => n8506, B2 => n9405, C1 => n8331, C2 => 
                           n9402, A => n1574, ZN => n1569);
   U848 : OAI221_X1 port map( B1 => n8467, B2 => n9417, C1 => n8435, C2 => 
                           n9414, A => n1573, ZN => n1570);
   U849 : NOR4_X1 port map( A1 => n1550, A2 => n1551, A3 => n1552, A4 => n1553,
                           ZN => n1549);
   U850 : OAI221_X1 port map( B1 => n8595, B2 => n9393, C1 => n8324, C2 => 
                           n9390, A => n1557, ZN => n1550);
   U851 : OAI221_X1 port map( B1 => n8507, B2 => n9405, C1 => n8332, C2 => 
                           n9402, A => n1556, ZN => n1551);
   U852 : OAI221_X1 port map( B1 => n8468, B2 => n9417, C1 => n8436, C2 => 
                           n9414, A => n1555, ZN => n1552);
   U853 : NOR4_X1 port map( A1 => n1532, A2 => n1533, A3 => n1534, A4 => n1535,
                           ZN => n1531);
   U854 : OAI221_X1 port map( B1 => n8596, B2 => n9393, C1 => n8325, C2 => 
                           n9390, A => n1539, ZN => n1532);
   U855 : OAI221_X1 port map( B1 => n8508, B2 => n9405, C1 => n8333, C2 => 
                           n9402, A => n1538, ZN => n1533);
   U856 : OAI221_X1 port map( B1 => n8469, B2 => n9417, C1 => n8437, C2 => 
                           n9414, A => n1537, ZN => n1534);
   U857 : NOR4_X1 port map( A1 => n1482, A2 => n1483, A3 => n1484, A4 => n1485,
                           ZN => n1481);
   U858 : OAI221_X1 port map( B1 => n8597, B2 => n9393, C1 => n8326, C2 => 
                           n9390, A => n1503, ZN => n1482);
   U859 : OAI221_X1 port map( B1 => n8509, B2 => n9405, C1 => n8334, C2 => 
                           n9402, A => n1498, ZN => n1483);
   U860 : OAI221_X1 port map( B1 => n8470, B2 => n9417, C1 => n8438, C2 => 
                           n9414, A => n1493, ZN => n1484);
   U861 : NOR4_X1 port map( A1 => n2090, A2 => n2091, A3 => n2092, A4 => n2093,
                           ZN => n2070);
   U862 : OAI221_X1 port map( B1 => n8886, B2 => n9343, C1 => n8862, C2 => 
                           n9340, A => n2099, ZN => n2090);
   U863 : OAI221_X1 port map( B1 => n8742, B2 => n9367, C1 => n8718, C2 => 
                           n9364, A => n2096, ZN => n2092);
   U864 : OAI221_X1 port map( B1 => n8798, B2 => n9355, C1 => n8774, C2 => 
                           n9352, A => n2097, ZN => n2091);
   U865 : NOR4_X1 port map( A1 => n2062, A2 => n2063, A3 => n2064, A4 => n2065,
                           ZN => n2052);
   U866 : OAI221_X1 port map( B1 => n8887, B2 => n9343, C1 => n8863, C2 => 
                           n9340, A => n2069, ZN => n2062);
   U867 : OAI221_X1 port map( B1 => n8743, B2 => n9367, C1 => n8719, C2 => 
                           n9364, A => n2067, ZN => n2064);
   U868 : OAI221_X1 port map( B1 => n8799, B2 => n9355, C1 => n8775, C2 => 
                           n9352, A => n2068, ZN => n2063);
   U869 : NOR4_X1 port map( A1 => n2044, A2 => n2045, A3 => n2046, A4 => n2047,
                           ZN => n2034);
   U870 : OAI221_X1 port map( B1 => n8888, B2 => n9343, C1 => n8864, C2 => 
                           n9340, A => n2051, ZN => n2044);
   U871 : OAI221_X1 port map( B1 => n8744, B2 => n9367, C1 => n8720, C2 => 
                           n9364, A => n2049, ZN => n2046);
   U872 : OAI221_X1 port map( B1 => n8800, B2 => n9355, C1 => n8776, C2 => 
                           n9352, A => n2050, ZN => n2045);
   U873 : NOR4_X1 port map( A1 => n2026, A2 => n2027, A3 => n2028, A4 => n2029,
                           ZN => n2016);
   U874 : OAI221_X1 port map( B1 => n8889, B2 => n9343, C1 => n8865, C2 => 
                           n9340, A => n2033, ZN => n2026);
   U875 : OAI221_X1 port map( B1 => n8745, B2 => n9367, C1 => n8721, C2 => 
                           n9364, A => n2031, ZN => n2028);
   U876 : OAI221_X1 port map( B1 => n8801, B2 => n9355, C1 => n8777, C2 => 
                           n9352, A => n2032, ZN => n2027);
   U877 : NOR4_X1 port map( A1 => n2008, A2 => n2009, A3 => n2010, A4 => n2011,
                           ZN => n1998);
   U878 : OAI221_X1 port map( B1 => n8890, B2 => n9343, C1 => n8866, C2 => 
                           n9340, A => n2015, ZN => n2008);
   U879 : OAI221_X1 port map( B1 => n8746, B2 => n9367, C1 => n8722, C2 => 
                           n9364, A => n2013, ZN => n2010);
   U880 : OAI221_X1 port map( B1 => n8802, B2 => n9355, C1 => n8778, C2 => 
                           n9352, A => n2014, ZN => n2009);
   U881 : NOR4_X1 port map( A1 => n1990, A2 => n1991, A3 => n1992, A4 => n1993,
                           ZN => n1980);
   U882 : OAI221_X1 port map( B1 => n8891, B2 => n9343, C1 => n8867, C2 => 
                           n9340, A => n1997, ZN => n1990);
   U883 : OAI221_X1 port map( B1 => n8747, B2 => n9367, C1 => n8723, C2 => 
                           n9364, A => n1995, ZN => n1992);
   U884 : OAI221_X1 port map( B1 => n8803, B2 => n9355, C1 => n8779, C2 => 
                           n9352, A => n1996, ZN => n1991);
   U885 : NOR4_X1 port map( A1 => n1972, A2 => n1973, A3 => n1974, A4 => n1975,
                           ZN => n1962);
   U886 : OAI221_X1 port map( B1 => n8892, B2 => n9343, C1 => n8868, C2 => 
                           n9340, A => n1979, ZN => n1972);
   U887 : OAI221_X1 port map( B1 => n8748, B2 => n9367, C1 => n8724, C2 => 
                           n9364, A => n1977, ZN => n1974);
   U888 : OAI221_X1 port map( B1 => n8804, B2 => n9355, C1 => n8780, C2 => 
                           n9352, A => n1978, ZN => n1973);
   U889 : NOR4_X1 port map( A1 => n1954, A2 => n1955, A3 => n1956, A4 => n1957,
                           ZN => n1944);
   U890 : OAI221_X1 port map( B1 => n8893, B2 => n9343, C1 => n8869, C2 => 
                           n9340, A => n1961, ZN => n1954);
   U891 : OAI221_X1 port map( B1 => n8749, B2 => n9367, C1 => n8725, C2 => 
                           n9364, A => n1959, ZN => n1956);
   U892 : OAI221_X1 port map( B1 => n8805, B2 => n9355, C1 => n8781, C2 => 
                           n9352, A => n1960, ZN => n1955);
   U893 : NAND2_X1 port map( A1 => n982, A2 => n983, ZN => OUT1(26));
   U894 : NOR4_X1 port map( A1 => n984, A2 => n985, A3 => n986, A4 => n987, ZN 
                           => n983);
   U895 : NOR4_X1 port map( A1 => n992, A2 => n993, A3 => n994, A4 => n995, ZN 
                           => n982);
   U896 : OAI221_X1 port map( B1 => n2143, B2 => n9489, C1 => n8401, C2 => 
                           n9486, A => n991, ZN => n984);
   U897 : AND3_X1 port map( A1 => n849, A2 => n9918, A3 => ADD_WR(4), ZN => 
                           n816);
   U898 : AND3_X1 port map( A1 => ADD_WR(4), A2 => n849, A3 => ADD_WR(3), ZN =>
                           n821);
   U899 : AND3_X1 port map( A1 => n849, A2 => n9917, A3 => ADD_WR(3), ZN => 
                           n826);
   U900 : OAI221_X1 port map( B1 => n8658, B2 => n9475, C1 => n8634, C2 => 
                           n9472, A => n1392, ZN => n1391);
   U901 : AOI22_X1 port map( A1 => n9469, A2 => n10189, B1 => n9468, B2 => 
                           n10253, ZN => n1392);
   U902 : OAI221_X1 port map( B1 => n8659, B2 => n9475, C1 => n8635, C2 => 
                           n9472, A => n1374, ZN => n1373);
   U903 : AOI22_X1 port map( A1 => n9469, A2 => n10188, B1 => n9468, B2 => 
                           n10252, ZN => n1374);
   U904 : OAI221_X1 port map( B1 => n8674, B2 => n9476, C1 => n8650, C2 => 
                           n9473, A => n1104, ZN => n1103);
   U905 : AOI22_X1 port map( A1 => n9470, A2 => n10173, B1 => n9466, B2 => 
                           n10237, ZN => n1104);
   U906 : OAI221_X1 port map( B1 => n8669, B2 => n9476, C1 => n8645, C2 => 
                           n9473, A => n1194, ZN => n1193);
   U907 : AOI22_X1 port map( A1 => n9470, A2 => n10178, B1 => n9467, B2 => 
                           n10242, ZN => n1194);
   U908 : OAI221_X1 port map( B1 => n8675, B2 => n9476, C1 => n8651, C2 => 
                           n9473, A => n1086, ZN => n1085);
   U909 : AOI22_X1 port map( A1 => n9470, A2 => n10172, B1 => n9466, B2 => 
                           n10236, ZN => n1086);
   U910 : OAI221_X1 port map( B1 => n8665, B2 => n9475, C1 => n8641, C2 => 
                           n9472, A => n1266, ZN => n1265);
   U911 : AOI22_X1 port map( A1 => n9469, A2 => n10182, B1 => n9467, B2 => 
                           n10246, ZN => n1266);
   U912 : OAI221_X1 port map( B1 => n8676, B2 => n9476, C1 => n8652, C2 => 
                           n9473, A => n1068, ZN => n1067);
   U913 : AOI22_X1 port map( A1 => n9470, A2 => n10171, B1 => n9466, B2 => 
                           n10235, ZN => n1068);
   U914 : OAI221_X1 port map( B1 => n8670, B2 => n9476, C1 => n8646, C2 => 
                           n9473, A => n1176, ZN => n1175);
   U915 : AOI22_X1 port map( A1 => n9470, A2 => n10177, B1 => n9467, B2 => 
                           n10241, ZN => n1176);
   U916 : OAI221_X1 port map( B1 => n8666, B2 => n9476, C1 => n8642, C2 => 
                           n9473, A => n1248, ZN => n1247);
   U917 : AOI22_X1 port map( A1 => n9470, A2 => n10181, B1 => n9467, B2 => 
                           n10245, ZN => n1248);
   U918 : OAI221_X1 port map( B1 => n8677, B2 => n9476, C1 => n8653, C2 => 
                           n9473, A => n1050, ZN => n1049);
   U919 : AOI22_X1 port map( A1 => n9470, A2 => n10170, B1 => n9466, B2 => 
                           n10234, ZN => n1050);
   U920 : OAI221_X1 port map( B1 => n8673, B2 => n9476, C1 => n8649, C2 => 
                           n9473, A => n1122, ZN => n1121);
   U921 : AOI22_X1 port map( A1 => n9470, A2 => n10174, B1 => n9467, B2 => 
                           n10238, ZN => n1122);
   U922 : OAI221_X1 port map( B1 => n8655, B2 => n9475, C1 => n8631, C2 => 
                           n9472, A => n1446, ZN => n1445);
   U923 : AOI22_X1 port map( A1 => n9469, A2 => n10192, B1 => n9468, B2 => 
                           n10256, ZN => n1446);
   U924 : OAI221_X1 port map( B1 => n8679, B2 => n9477, C1 => n8296, C2 => 
                           n9474, A => n1014, ZN => n1013);
   U925 : AOI22_X1 port map( A1 => n9471, A2 => n10584, B1 => n9466, B2 => 
                           n10232, ZN => n1014);
   U926 : OAI221_X1 port map( B1 => n8656, B2 => n9475, C1 => n8632, C2 => 
                           n9472, A => n1428, ZN => n1427);
   U927 : AOI22_X1 port map( A1 => n9469, A2 => n10191, B1 => n9468, B2 => 
                           n10255, ZN => n1428);
   U928 : OAI221_X1 port map( B1 => n8661, B2 => n9475, C1 => n8637, C2 => 
                           n9472, A => n1338, ZN => n1337);
   U929 : AOI22_X1 port map( A1 => n9469, A2 => n10186, B1 => n9468, B2 => 
                           n10250, ZN => n1338);
   U930 : OAI221_X1 port map( B1 => n8680, B2 => n9477, C1 => n8297, C2 => 
                           n9474, A => n996, ZN => n995);
   U931 : AOI22_X1 port map( A1 => n9471, A2 => n10583, B1 => n9466, B2 => 
                           n10231, ZN => n996);
   U932 : OAI221_X1 port map( B1 => n8662, B2 => n9475, C1 => n8638, C2 => 
                           n9472, A => n1320, ZN => n1319);
   U933 : AOI22_X1 port map( A1 => n9469, A2 => n10185, B1 => n9467, B2 => 
                           n10249, ZN => n1320);
   U934 : OAI221_X1 port map( B1 => n8684, B2 => n9477, C1 => n8301, C2 => 
                           n9474, A => n924, ZN => n923);
   U935 : AOI22_X1 port map( A1 => n9471, A2 => n10579, B1 => n9466, B2 => 
                           n10227, ZN => n924);
   U936 : OAI221_X1 port map( B1 => n8681, B2 => n9477, C1 => n8298, C2 => 
                           n9474, A => n978, ZN => n977);
   U937 : AOI22_X1 port map( A1 => n9471, A2 => n10582, B1 => n9466, B2 => 
                           n10230, ZN => n978);
   U938 : OAI221_X1 port map( B1 => n8663, B2 => n9475, C1 => n8639, C2 => 
                           n9472, A => n1302, ZN => n1301);
   U939 : AOI22_X1 port map( A1 => n9469, A2 => n10184, B1 => n9467, B2 => 
                           n10248, ZN => n1302);
   U940 : OAI221_X1 port map( B1 => n8662, B2 => n9379, C1 => n8638, C2 => 
                           n9376, A => n1940, ZN => n1939);
   U941 : AOI22_X1 port map( A1 => n9373, A2 => n10217, B1 => n9371, B2 => 
                           n10249, ZN => n1940);
   U942 : OAI221_X1 port map( B1 => n8663, B2 => n9379, C1 => n8639, C2 => 
                           n9376, A => n1922, ZN => n1921);
   U943 : AOI22_X1 port map( A1 => n9373, A2 => n10216, B1 => n9371, B2 => 
                           n10248, ZN => n1922);
   U944 : OAI221_X1 port map( B1 => n8664, B2 => n9379, C1 => n8640, C2 => 
                           n9376, A => n1904, ZN => n1903);
   U945 : AOI22_X1 port map( A1 => n9373, A2 => n10215, B1 => n9371, B2 => 
                           n10247, ZN => n1904);
   U946 : OAI221_X1 port map( B1 => n8665, B2 => n9379, C1 => n8641, C2 => 
                           n9376, A => n1886, ZN => n1885);
   U947 : AOI22_X1 port map( A1 => n9373, A2 => n10214, B1 => n9371, B2 => 
                           n10246, ZN => n1886);
   U948 : OAI221_X1 port map( B1 => n8666, B2 => n9380, C1 => n8642, C2 => 
                           n9377, A => n1868, ZN => n1867);
   U949 : AOI22_X1 port map( A1 => n9374, A2 => n10213, B1 => n9371, B2 => 
                           n10245, ZN => n1868);
   U950 : OAI221_X1 port map( B1 => n8668, B2 => n9380, C1 => n8644, C2 => 
                           n9377, A => n1832, ZN => n1831);
   U951 : AOI22_X1 port map( A1 => n9374, A2 => n10211, B1 => n9371, B2 => 
                           n10243, ZN => n1832);
   U952 : OAI221_X1 port map( B1 => n8669, B2 => n9380, C1 => n8645, C2 => 
                           n9377, A => n1814, ZN => n1813);
   U953 : AOI22_X1 port map( A1 => n9374, A2 => n10210, B1 => n9371, B2 => 
                           n10242, ZN => n1814);
   U954 : OAI221_X1 port map( B1 => n8670, B2 => n9380, C1 => n8646, C2 => 
                           n9377, A => n1796, ZN => n1795);
   U955 : AOI22_X1 port map( A1 => n9374, A2 => n10209, B1 => n9371, B2 => 
                           n10241, ZN => n1796);
   U956 : OAI221_X1 port map( B1 => n8672, B2 => n9380, C1 => n8648, C2 => 
                           n9377, A => n1760, ZN => n1759);
   U957 : AOI22_X1 port map( A1 => n9374, A2 => n10207, B1 => n9371, B2 => 
                           n10239, ZN => n1760);
   U958 : OAI221_X1 port map( B1 => n8673, B2 => n9380, C1 => n8649, C2 => 
                           n9377, A => n1742, ZN => n1741);
   U959 : AOI22_X1 port map( A1 => n9374, A2 => n10206, B1 => n9371, B2 => 
                           n10238, ZN => n1742);
   U960 : OAI221_X1 port map( B1 => n8674, B2 => n9380, C1 => n8650, C2 => 
                           n9377, A => n1724, ZN => n1723);
   U961 : AOI22_X1 port map( A1 => n9374, A2 => n10205, B1 => n9370, B2 => 
                           n10237, ZN => n1724);
   U962 : OAI221_X1 port map( B1 => n8675, B2 => n9380, C1 => n8651, C2 => 
                           n9377, A => n1706, ZN => n1705);
   U963 : AOI22_X1 port map( A1 => n9374, A2 => n10204, B1 => n9370, B2 => 
                           n10236, ZN => n1706);
   U964 : OAI221_X1 port map( B1 => n8676, B2 => n9380, C1 => n8652, C2 => 
                           n9377, A => n1688, ZN => n1687);
   U965 : AOI22_X1 port map( A1 => n9374, A2 => n10203, B1 => n9370, B2 => 
                           n10235, ZN => n1688);
   U966 : OAI221_X1 port map( B1 => n8677, B2 => n9380, C1 => n8653, C2 => 
                           n9377, A => n1670, ZN => n1669);
   U967 : AOI22_X1 port map( A1 => n9374, A2 => n10202, B1 => n9370, B2 => 
                           n10234, ZN => n1670);
   U968 : OAI221_X1 port map( B1 => n8678, B2 => n9381, C1 => n8295, C2 => 
                           n9378, A => n1652, ZN => n1651);
   U969 : AOI22_X1 port map( A1 => n9375, A2 => n10201, B1 => n9370, B2 => 
                           n10233, ZN => n1652);
   U970 : OAI221_X1 port map( B1 => n8679, B2 => n9381, C1 => n8296, C2 => 
                           n9378, A => n1634, ZN => n1633);
   U971 : AOI22_X1 port map( A1 => n9375, A2 => n10200, B1 => n9370, B2 => 
                           n10232, ZN => n1634);
   U972 : OAI221_X1 port map( B1 => n8680, B2 => n9381, C1 => n8297, C2 => 
                           n9378, A => n1616, ZN => n1615);
   U973 : AOI22_X1 port map( A1 => n9375, A2 => n10199, B1 => n9370, B2 => 
                           n10231, ZN => n1616);
   U974 : OAI221_X1 port map( B1 => n8681, B2 => n9381, C1 => n8298, C2 => 
                           n9378, A => n1598, ZN => n1597);
   U975 : AOI22_X1 port map( A1 => n9375, A2 => n10198, B1 => n9370, B2 => 
                           n10230, ZN => n1598);
   U976 : OAI221_X1 port map( B1 => n8682, B2 => n9381, C1 => n8299, C2 => 
                           n9378, A => n1580, ZN => n1579);
   U977 : AOI22_X1 port map( A1 => n9375, A2 => n10197, B1 => n9370, B2 => 
                           n10229, ZN => n1580);
   U978 : OAI221_X1 port map( B1 => n8683, B2 => n9381, C1 => n8300, C2 => 
                           n9378, A => n1562, ZN => n1561);
   U979 : AOI22_X1 port map( A1 => n9375, A2 => n10196, B1 => n9370, B2 => 
                           n10228, ZN => n1562);
   U980 : OAI221_X1 port map( B1 => n8684, B2 => n9381, C1 => n8301, C2 => 
                           n9378, A => n1544, ZN => n1543);
   U981 : AOI22_X1 port map( A1 => n9375, A2 => n10195, B1 => n9370, B2 => 
                           n10227, ZN => n1544);
   U982 : OAI221_X1 port map( B1 => n8685, B2 => n9381, C1 => n8302, C2 => 
                           n9378, A => n1512, ZN => n1509);
   U983 : AOI22_X1 port map( A1 => n9375, A2 => n10194, B1 => n9370, B2 => 
                           n10226, ZN => n1512);
   U984 : OAI221_X1 port map( B1 => n8601, B2 => n9523, C1 => n8569, C2 => 
                           n9520, A => n1402, ZN => n1401);
   U985 : AOI22_X1 port map( A1 => n9517, A2 => n10470, B1 => n9516, B2 => 
                           n10286, ZN => n1402);
   U986 : OAI221_X1 port map( B1 => n8602, B2 => n9523, C1 => n8570, C2 => 
                           n9520, A => n1384, ZN => n1383);
   U987 : AOI22_X1 port map( A1 => n9517, A2 => n10469, B1 => n9516, B2 => 
                           n10285, ZN => n1384);
   U988 : OAI221_X1 port map( B1 => n8603, B2 => n9523, C1 => n8571, C2 => 
                           n9520, A => n1366, ZN => n1365);
   U989 : AOI22_X1 port map( A1 => n9517, A2 => n10468, B1 => n9516, B2 => 
                           n10284, ZN => n1366);
   U990 : OAI221_X1 port map( B1 => n8618, B2 => n9524, C1 => n8586, C2 => 
                           n9521, A => n1096, ZN => n1095);
   U991 : AOI22_X1 port map( A1 => n9518, A2 => n10453, B1 => n9514, B2 => 
                           n10269, ZN => n1096);
   U992 : OAI221_X1 port map( B1 => n8608, B2 => n9523, C1 => n8576, C2 => 
                           n9520, A => n1276, ZN => n1275);
   U993 : AOI22_X1 port map( A1 => n9517, A2 => n10463, B1 => n9515, B2 => 
                           n10279, ZN => n1276);
   U994 : OAI221_X1 port map( B1 => n8609, B2 => n9523, C1 => n8577, C2 => 
                           n9520, A => n1258, ZN => n1257);
   U995 : AOI22_X1 port map( A1 => n9517, A2 => n10462, B1 => n9515, B2 => 
                           n10278, ZN => n1258);
   U996 : OAI221_X1 port map( B1 => n8620, B2 => n9524, C1 => n8588, C2 => 
                           n9521, A => n1060, ZN => n1059);
   U997 : AOI22_X1 port map( A1 => n9518, A2 => n10451, B1 => n9514, B2 => 
                           n10267, ZN => n1060);
   U998 : OAI221_X1 port map( B1 => n8619, B2 => n9524, C1 => n8587, C2 => 
                           n9521, A => n1078, ZN => n1077);
   U999 : AOI22_X1 port map( A1 => n9518, A2 => n10452, B1 => n9514, B2 => 
                           n10268, ZN => n1078);
   U1000 : OAI221_X1 port map( B1 => n8614, B2 => n9524, C1 => n8582, C2 => 
                           n9521, A => n1168, ZN => n1167);
   U1001 : AOI22_X1 port map( A1 => n9518, A2 => n10457, B1 => n9515, B2 => 
                           n10273, ZN => n1168);
   U1002 : OAI221_X1 port map( B1 => n8610, B2 => n9524, C1 => n8578, C2 => 
                           n9521, A => n1240, ZN => n1239);
   U1003 : AOI22_X1 port map( A1 => n9518, A2 => n10461, B1 => n9515, B2 => 
                           n10277, ZN => n1240);
   U1004 : OAI221_X1 port map( B1 => n8621, B2 => n9524, C1 => n8589, C2 => 
                           n9521, A => n1042, ZN => n1041);
   U1005 : AOI22_X1 port map( A1 => n9518, A2 => n10450, B1 => n9514, B2 => 
                           n10266, ZN => n1042);
   U1006 : OAI221_X1 port map( B1 => n8599, B2 => n9523, C1 => n8567, C2 => 
                           n9520, A => n1438, ZN => n1437);
   U1007 : AOI22_X1 port map( A1 => n9517, A2 => n10472, B1 => n9516, B2 => 
                           n10288, ZN => n1438);
   U1008 : OAI221_X1 port map( B1 => n8600, B2 => n9523, C1 => n8568, C2 => 
                           n9520, A => n1420, ZN => n1419);
   U1009 : AOI22_X1 port map( A1 => n9517, A2 => n10471, B1 => n9516, B2 => 
                           n10287, ZN => n1420);
   U1010 : OAI221_X1 port map( B1 => n8604, B2 => n9523, C1 => n8572, C2 => 
                           n9520, A => n1348, ZN => n1347);
   U1011 : AOI22_X1 port map( A1 => n9517, A2 => n10467, B1 => n9516, B2 => 
                           n10283, ZN => n1348);
   U1012 : OAI221_X1 port map( B1 => n8622, B2 => n9525, C1 => n8590, C2 => 
                           n9522, A => n1024, ZN => n1023);
   U1013 : AOI22_X1 port map( A1 => n9519, A2 => n10449, B1 => n9514, B2 => 
                           n10265, ZN => n1024);
   U1014 : OAI221_X1 port map( B1 => n8627, B2 => n9525, C1 => n8595, C2 => 
                           n9522, A => n934, ZN => n933);
   U1015 : AOI22_X1 port map( A1 => n9519, A2 => n10444, B1 => n9514, B2 => 
                           n10260, ZN => n934);
   U1016 : OAI221_X1 port map( B1 => n8605, B2 => n9523, C1 => n8573, C2 => 
                           n9520, A => n1330, ZN => n1329);
   U1017 : AOI22_X1 port map( A1 => n9517, A2 => n10466, B1 => n9516, B2 => 
                           n10282, ZN => n1330);
   U1018 : OAI221_X1 port map( B1 => n8624, B2 => n9525, C1 => n8592, C2 => 
                           n9522, A => n988, ZN => n987);
   U1019 : AOI22_X1 port map( A1 => n9519, A2 => n10447, B1 => n9514, B2 => 
                           n10263, ZN => n988);
   U1020 : OAI221_X1 port map( B1 => n8628, B2 => n9525, C1 => n8596, C2 => 
                           n9522, A => n916, ZN => n915);
   U1021 : AOI22_X1 port map( A1 => n9519, A2 => n10443, B1 => n9514, B2 => 
                           n10259, ZN => n916);
   U1022 : OAI221_X1 port map( B1 => n8606, B2 => n9523, C1 => n8574, C2 => 
                           n9520, A => n1312, ZN => n1311);
   U1023 : AOI22_X1 port map( A1 => n9517, A2 => n10465, B1 => n9515, B2 => 
                           n10281, ZN => n1312);
   U1024 : OAI221_X1 port map( B1 => n8625, B2 => n9525, C1 => n8593, C2 => 
                           n9522, A => n970, ZN => n969);
   U1025 : AOI22_X1 port map( A1 => n9519, A2 => n10446, B1 => n9514, B2 => 
                           n10262, ZN => n970);
   U1026 : OAI221_X1 port map( B1 => n8607, B2 => n9523, C1 => n8575, C2 => 
                           n9520, A => n1294, ZN => n1293);
   U1027 : AOI22_X1 port map( A1 => n9517, A2 => n10464, B1 => n9515, B2 => 
                           n10280, ZN => n1294);
   U1028 : OAI221_X1 port map( B1 => n8667, B2 => n9380, C1 => n8643, C2 => 
                           n9377, A => n1850, ZN => n1849);
   U1029 : AOI22_X1 port map( A1 => n9374, A2 => n10212, B1 => n9371, B2 => 
                           n10244, ZN => n1850);
   U1030 : OAI221_X1 port map( B1 => n8671, B2 => n9380, C1 => n8647, C2 => 
                           n9377, A => n1778, ZN => n1777);
   U1031 : AOI22_X1 port map( A1 => n9374, A2 => n10208, B1 => n9371, B2 => 
                           n10240, ZN => n1778);
   U1032 : OAI221_X1 port map( B1 => n8778, B2 => n9463, C1 => n8237, C2 => 
                           n9460, A => n1393, ZN => n1390);
   U1033 : AOI22_X1 port map( A1 => n9457, A2 => n10133, B1 => n9456, B2 => 
                           n10165, ZN => n1393);
   U1034 : OAI221_X1 port map( B1 => n8334, B2 => n9513, C1 => n8182, C2 => 
                           n9510, A => n873, ZN => n864);
   U1035 : AOI22_X1 port map( A1 => n9507, A2 => n10538, B1 => n9502, B2 => 
                           n10410, ZN => n873);
   U1036 : OAI221_X1 port map( B1 => n8779, B2 => n9463, C1 => n8235, C2 => 
                           n9460, A => n1375, ZN => n1372);
   U1037 : AOI22_X1 port map( A1 => n9457, A2 => n10132, B1 => n9456, B2 => 
                           n10164, ZN => n1375);
   U1038 : OAI221_X1 port map( B1 => n8794, B2 => n9464, C1 => n8205, C2 => 
                           n9461, A => n1105, ZN => n1102);
   U1039 : AOI22_X1 port map( A1 => n9458, A2 => n10117, B1 => n9454, B2 => 
                           n10149, ZN => n1105);
   U1040 : OAI221_X1 port map( B1 => n8789, B2 => n9464, C1 => n8215, C2 => 
                           n9461, A => n1195, ZN => n1192);
   U1041 : AOI22_X1 port map( A1 => n9458, A2 => n10122, B1 => n9455, B2 => 
                           n10154, ZN => n1195);
   U1042 : OAI221_X1 port map( B1 => n8795, B2 => n9464, C1 => n8203, C2 => 
                           n9461, A => n1087, ZN => n1084);
   U1043 : AOI22_X1 port map( A1 => n9458, A2 => n10116, B1 => n9454, B2 => 
                           n10148, ZN => n1087);
   U1044 : OAI221_X1 port map( B1 => n8785, B2 => n9463, C1 => n8223, C2 => 
                           n9460, A => n1267, ZN => n1264);
   U1045 : AOI22_X1 port map( A1 => n9457, A2 => n10126, B1 => n9455, B2 => 
                           n10158, ZN => n1267);
   U1046 : OAI221_X1 port map( B1 => n8796, B2 => n9464, C1 => n8201, C2 => 
                           n9461, A => n1069, ZN => n1066);
   U1047 : AOI22_X1 port map( A1 => n9458, A2 => n10115, B1 => n9454, B2 => 
                           n10147, ZN => n1069);
   U1048 : OAI221_X1 port map( B1 => n8471, B2 => n9511, C1 => n8244, C2 => 
                           n9508, A => n1462, ZN => n1454);
   U1049 : AOI22_X1 port map( A1 => n9505, A2 => n10609, B1 => n9504, B2 => 
                           n10441, ZN => n1462);
   U1050 : OAI221_X1 port map( B1 => n8790, B2 => n9464, C1 => n8213, C2 => 
                           n9461, A => n1177, ZN => n1174);
   U1051 : AOI22_X1 port map( A1 => n9458, A2 => n10121, B1 => n9455, B2 => 
                           n10153, ZN => n1177);
   U1052 : OAI221_X1 port map( B1 => n8786, B2 => n9464, C1 => n8221, C2 => 
                           n9461, A => n1249, ZN => n1246);
   U1053 : AOI22_X1 port map( A1 => n9458, A2 => n10125, B1 => n9455, B2 => 
                           n10157, ZN => n1249);
   U1054 : OAI221_X1 port map( B1 => n8797, B2 => n9464, C1 => n8199, C2 => 
                           n9461, A => n1051, ZN => n1048);
   U1055 : AOI22_X1 port map( A1 => n9458, A2 => n10114, B1 => n9454, B2 => 
                           n10146, ZN => n1051);
   U1056 : OAI221_X1 port map( B1 => n8793, B2 => n9464, C1 => n8207, C2 => 
                           n9461, A => n1123, ZN => n1120);
   U1057 : AOI22_X1 port map( A1 => n9458, A2 => n10118, B1 => n9455, B2 => 
                           n10150, ZN => n1123);
   U1058 : OAI221_X1 port map( B1 => n8775, B2 => n9463, C1 => n8243, C2 => 
                           n9460, A => n1447, ZN => n1444);
   U1059 : AOI22_X1 port map( A1 => n9457, A2 => n10136, B1 => n9456, B2 => 
                           n10168, ZN => n1447);
   U1060 : OAI221_X1 port map( B1 => n8312, B2 => n9465, C1 => n8195, C2 => 
                           n9462, A => n1015, ZN => n1012);
   U1061 : AOI22_X1 port map( A1 => n9459, A2 => n10112, B1 => n9454, B2 => 
                           n10144, ZN => n1015);
   U1062 : OAI221_X1 port map( B1 => n8776, B2 => n9463, C1 => n8241, C2 => 
                           n9460, A => n1429, ZN => n1426);
   U1063 : AOI22_X1 port map( A1 => n9457, A2 => n10135, B1 => n9456, B2 => 
                           n10167, ZN => n1429);
   U1064 : OAI221_X1 port map( B1 => n8781, B2 => n9463, C1 => n8231, C2 => 
                           n9460, A => n1339, ZN => n1336);
   U1065 : AOI22_X1 port map( A1 => n9457, A2 => n10130, B1 => n9456, B2 => 
                           n10162, ZN => n1339);
   U1066 : OAI221_X1 port map( B1 => n8313, B2 => n9465, C1 => n8193, C2 => 
                           n9462, A => n997, ZN => n994);
   U1067 : AOI22_X1 port map( A1 => n9459, A2 => n10111, B1 => n9454, B2 => 
                           n10143, ZN => n997);
   U1068 : OAI221_X1 port map( B1 => n8328, B2 => n9513, C1 => n8194, C2 => 
                           n9510, A => n1007, ZN => n1004);
   U1069 : AOI22_X1 port map( A1 => n9507, A2 => n10544, B1 => n9502, B2 => 
                           n10416, ZN => n1007);
   U1070 : OAI221_X1 port map( B1 => n8331, B2 => n9513, C1 => n8188, C2 => 
                           n9510, A => n953, ZN => n950);
   U1071 : AOI22_X1 port map( A1 => n9507, A2 => n10541, B1 => n9502, B2 => 
                           n10413, ZN => n953);
   U1072 : OAI221_X1 port map( B1 => n8327, B2 => n9513, C1 => n8196, C2 => 
                           n9510, A => n1025, ZN => n1022);
   U1073 : AOI22_X1 port map( A1 => n9507, A2 => n10545, B1 => n9502, B2 => 
                           n10417, ZN => n1025);
   U1074 : OAI221_X1 port map( B1 => n8332, B2 => n9513, C1 => n8186, C2 => 
                           n9510, A => n935, ZN => n932);
   U1075 : AOI22_X1 port map( A1 => n9507, A2 => n10540, B1 => n9502, B2 => 
                           n10412, ZN => n935);
   U1076 : OAI221_X1 port map( B1 => n8782, B2 => n9463, C1 => n8229, C2 => 
                           n9460, A => n1321, ZN => n1318);
   U1077 : AOI22_X1 port map( A1 => n9457, A2 => n10129, B1 => n9455, B2 => 
                           n10161, ZN => n1321);
   U1078 : OAI221_X1 port map( B1 => n8317, B2 => n9465, C1 => n8185, C2 => 
                           n9462, A => n925, ZN => n922);
   U1079 : AOI22_X1 port map( A1 => n9459, A2 => n10107, B1 => n9454, B2 => 
                           n10139, ZN => n925);
   U1080 : OAI221_X1 port map( B1 => n8329, B2 => n9513, C1 => n8192, C2 => 
                           n9510, A => n989, ZN => n986);
   U1081 : AOI22_X1 port map( A1 => n9507, A2 => n10543, B1 => n9502, B2 => 
                           n10415, ZN => n989);
   U1082 : OAI221_X1 port map( B1 => n8314, B2 => n9465, C1 => n8191, C2 => 
                           n9462, A => n979, ZN => n976);
   U1083 : AOI22_X1 port map( A1 => n9459, A2 => n10110, B1 => n9454, B2 => 
                           n10142, ZN => n979);
   U1084 : OAI221_X1 port map( B1 => n8783, B2 => n9463, C1 => n8227, C2 => 
                           n9460, A => n1303, ZN => n1300);
   U1085 : AOI22_X1 port map( A1 => n9457, A2 => n10128, B1 => n9455, B2 => 
                           n10160, ZN => n1303);
   U1086 : OAI221_X1 port map( B1 => n8477, B2 => n9511, C1 => n8232, C2 => 
                           n9508, A => n1349, ZN => n1346);
   U1087 : AOI22_X1 port map( A1 => n9505, A2 => n10603, B1 => n9504, B2 => 
                           n10435, ZN => n1349);
   U1088 : OAI221_X1 port map( B1 => n8333, B2 => n9513, C1 => n8184, C2 => 
                           n9510, A => n917, ZN => n914);
   U1089 : AOI22_X1 port map( A1 => n9507, A2 => n10539, B1 => n9502, B2 => 
                           n10411, ZN => n917);
   U1090 : OAI221_X1 port map( B1 => n8330, B2 => n9513, C1 => n8190, C2 => 
                           n9510, A => n971, ZN => n968);
   U1091 : AOI22_X1 port map( A1 => n9507, A2 => n10542, B1 => n9502, B2 => 
                           n10414, ZN => n971);
   U1092 : OAI221_X1 port map( B1 => n8513, B2 => n9499, C1 => n8481, C2 => 
                           n9496, A => n1404, ZN => n1399);
   U1093 : AOI22_X1 port map( A1 => n9493, A2 => n10502, B1 => n9492, B2 => 
                           n10374, ZN => n1404);
   U1094 : OAI221_X1 port map( B1 => n8541, B2 => n9501, C1 => n8509, C2 => 
                           n9498, A => n878, ZN => n863);
   U1095 : AOI22_X1 port map( A1 => n9495, A2 => n10474, B1 => n9490, B2 => 
                           n10346, ZN => n878);
   U1096 : OAI221_X1 port map( B1 => n8514, B2 => n9499, C1 => n8482, C2 => 
                           n9496, A => n1386, ZN => n1381);
   U1097 : AOI22_X1 port map( A1 => n9493, A2 => n10501, B1 => n9492, B2 => 
                           n10373, ZN => n1386);
   U1098 : OAI221_X1 port map( B1 => n8834, B2 => n9451, C1 => n8802, C2 => 
                           n9448, A => n1394, ZN => n1389);
   U1099 : AOI22_X1 port map( A1 => n9445, A2 => n10005, B1 => n9444, B2 => 
                           n10037, ZN => n1394);
   U1100 : OAI221_X1 port map( B1 => n8515, B2 => n9499, C1 => n8483, C2 => 
                           n9496, A => n1368, ZN => n1363);
   U1101 : AOI22_X1 port map( A1 => n9493, A2 => n10500, B1 => n9492, B2 => 
                           n10372, ZN => n1368);
   U1102 : OAI221_X1 port map( B1 => n8835, B2 => n9451, C1 => n8803, C2 => 
                           n9448, A => n1376, ZN => n1371);
   U1103 : AOI22_X1 port map( A1 => n9445, A2 => n10004, B1 => n9444, B2 => 
                           n10036, ZN => n1376);
   U1104 : OAI221_X1 port map( B1 => n8523, B2 => n9500, C1 => n8491, C2 => 
                           n9497, A => n1224, ZN => n1219);
   U1105 : AOI22_X1 port map( A1 => n9494, A2 => n10492, B1 => n9491, B2 => 
                           n10364, ZN => n1224);
   U1106 : OAI221_X1 port map( B1 => n8510, B2 => n9499, C1 => n8478, C2 => 
                           n9496, A => n1465, ZN => n1453);
   U1107 : AOI22_X1 port map( A1 => n9493, A2 => n10505, B1 => n9492, B2 => 
                           n10377, ZN => n1465);
   U1108 : OAI221_X1 port map( B1 => n8524, B2 => n9500, C1 => n8492, C2 => 
                           n9497, A => n1206, ZN => n1201);
   U1109 : AOI22_X1 port map( A1 => n9494, A2 => n10491, B1 => n9491, B2 => 
                           n10363, ZN => n1206);
   U1110 : OAI221_X1 port map( B1 => n8525, B2 => n9500, C1 => n8493, C2 => 
                           n9497, A => n1188, ZN => n1183);
   U1111 : AOI22_X1 port map( A1 => n9494, A2 => n10490, B1 => n9491, B2 => 
                           n10362, ZN => n1188);
   U1112 : OAI221_X1 port map( B1 => n8530, B2 => n9500, C1 => n8498, C2 => 
                           n9497, A => n1098, ZN => n1093);
   U1113 : AOI22_X1 port map( A1 => n9494, A2 => n10485, B1 => n9490, B2 => 
                           n10357, ZN => n1098);
   U1114 : OAI221_X1 port map( B1 => n8850, B2 => n9452, C1 => n8818, C2 => 
                           n9449, A => n1106, ZN => n1101);
   U1115 : AOI22_X1 port map( A1 => n9446, A2 => n9989, B1 => n9442, B2 => 
                           n10021, ZN => n1106);
   U1116 : OAI221_X1 port map( B1 => n8845, B2 => n9452, C1 => n8813, C2 => 
                           n9449, A => n1196, ZN => n1191);
   U1117 : AOI22_X1 port map( A1 => n9446, A2 => n9994, B1 => n9443, B2 => 
                           n10026, ZN => n1196);
   U1118 : OAI221_X1 port map( B1 => n8520, B2 => n9499, C1 => n8488, C2 => 
                           n9496, A => n1278, ZN => n1273);
   U1119 : AOI22_X1 port map( A1 => n9493, A2 => n10495, B1 => n9491, B2 => 
                           n10367, ZN => n1278);
   U1120 : OAI221_X1 port map( B1 => n8521, B2 => n9499, C1 => n8489, C2 => 
                           n9496, A => n1260, ZN => n1255);
   U1121 : AOI22_X1 port map( A1 => n9493, A2 => n10494, B1 => n9491, B2 => 
                           n10366, ZN => n1260);
   U1122 : OAI221_X1 port map( B1 => n8532, B2 => n9500, C1 => n8500, C2 => 
                           n9497, A => n1062, ZN => n1057);
   U1123 : AOI22_X1 port map( A1 => n9494, A2 => n10483, B1 => n9490, B2 => 
                           n10355, ZN => n1062);
   U1124 : OAI221_X1 port map( B1 => n8531, B2 => n9500, C1 => n8499, C2 => 
                           n9497, A => n1080, ZN => n1075);
   U1125 : AOI22_X1 port map( A1 => n9494, A2 => n10484, B1 => n9490, B2 => 
                           n10356, ZN => n1080);
   U1126 : OAI221_X1 port map( B1 => n8851, B2 => n9452, C1 => n8819, C2 => 
                           n9449, A => n1088, ZN => n1083);
   U1127 : AOI22_X1 port map( A1 => n9446, A2 => n9988, B1 => n9442, B2 => 
                           n10020, ZN => n1088);
   U1128 : OAI221_X1 port map( B1 => n8841, B2 => n9451, C1 => n8809, C2 => 
                           n9448, A => n1268, ZN => n1263);
   U1129 : AOI22_X1 port map( A1 => n9445, A2 => n9998, B1 => n9443, B2 => 
                           n10030, ZN => n1268);
   U1130 : OAI221_X1 port map( B1 => n8852, B2 => n9452, C1 => n8820, C2 => 
                           n9449, A => n1070, ZN => n1065);
   U1131 : AOI22_X1 port map( A1 => n9446, A2 => n9987, B1 => n9442, B2 => 
                           n10019, ZN => n1070);
   U1132 : OAI221_X1 port map( B1 => n8526, B2 => n9500, C1 => n8494, C2 => 
                           n9497, A => n1170, ZN => n1165);
   U1133 : AOI22_X1 port map( A1 => n9494, A2 => n10489, B1 => n9491, B2 => 
                           n10361, ZN => n1170);
   U1134 : OAI221_X1 port map( B1 => n8846, B2 => n9452, C1 => n8814, C2 => 
                           n9449, A => n1178, ZN => n1173);
   U1135 : AOI22_X1 port map( A1 => n9446, A2 => n9993, B1 => n9443, B2 => 
                           n10025, ZN => n1178);
   U1136 : OAI221_X1 port map( B1 => n8522, B2 => n9500, C1 => n8490, C2 => 
                           n9497, A => n1242, ZN => n1237);
   U1137 : AOI22_X1 port map( A1 => n9494, A2 => n10493, B1 => n9491, B2 => 
                           n10365, ZN => n1242);
   U1138 : OAI221_X1 port map( B1 => n8533, B2 => n9500, C1 => n8501, C2 => 
                           n9497, A => n1044, ZN => n1039);
   U1139 : AOI22_X1 port map( A1 => n9494, A2 => n10482, B1 => n9490, B2 => 
                           n10354, ZN => n1044);
   U1140 : OAI221_X1 port map( B1 => n8842, B2 => n9452, C1 => n8810, C2 => 
                           n9449, A => n1250, ZN => n1245);
   U1141 : AOI22_X1 port map( A1 => n9446, A2 => n9997, B1 => n9443, B2 => 
                           n10029, ZN => n1250);
   U1142 : OAI221_X1 port map( B1 => n8853, B2 => n9452, C1 => n8821, C2 => 
                           n9449, A => n1052, ZN => n1047);
   U1143 : AOI22_X1 port map( A1 => n9446, A2 => n9986, B1 => n9442, B2 => 
                           n10018, ZN => n1052);
   U1144 : OAI221_X1 port map( B1 => n8527, B2 => n9500, C1 => n8495, C2 => 
                           n9497, A => n1152, ZN => n1147);
   U1145 : AOI22_X1 port map( A1 => n9494, A2 => n10488, B1 => n9491, B2 => 
                           n10360, ZN => n1152);
   U1146 : OAI221_X1 port map( B1 => n8528, B2 => n9500, C1 => n8496, C2 => 
                           n9497, A => n1134, ZN => n1129);
   U1147 : AOI22_X1 port map( A1 => n9494, A2 => n10487, B1 => n9491, B2 => 
                           n10359, ZN => n1134);
   U1148 : OAI221_X1 port map( B1 => n8529, B2 => n9500, C1 => n8497, C2 => 
                           n9497, A => n1116, ZN => n1111);
   U1149 : AOI22_X1 port map( A1 => n9494, A2 => n10486, B1 => n9491, B2 => 
                           n10358, ZN => n1116);
   U1150 : OAI221_X1 port map( B1 => n8849, B2 => n9452, C1 => n8817, C2 => 
                           n9449, A => n1124, ZN => n1119);
   U1151 : AOI22_X1 port map( A1 => n9446, A2 => n9990, B1 => n9443, B2 => 
                           n10022, ZN => n1124);
   U1152 : OAI221_X1 port map( B1 => n8511, B2 => n9499, C1 => n8479, C2 => 
                           n9496, A => n1440, ZN => n1435);
   U1153 : AOI22_X1 port map( A1 => n9493, A2 => n10504, B1 => n9492, B2 => 
                           n10376, ZN => n1440);
   U1154 : OAI221_X1 port map( B1 => n8831, B2 => n9451, C1 => n8799, C2 => 
                           n9448, A => n1448, ZN => n1443);
   U1155 : AOI22_X1 port map( A1 => n9445, A2 => n10008, B1 => n9444, B2 => 
                           n10040, ZN => n1448);
   U1156 : OAI221_X1 port map( B1 => n8512, B2 => n9499, C1 => n8480, C2 => 
                           n9496, A => n1422, ZN => n1417);
   U1157 : AOI22_X1 port map( A1 => n9493, A2 => n10503, B1 => n9492, B2 => 
                           n10375, ZN => n1422);
   U1158 : OAI221_X1 port map( B1 => n8535, B2 => n9501, C1 => n8503, C2 => 
                           n9498, A => n1008, ZN => n1003);
   U1159 : AOI22_X1 port map( A1 => n9495, A2 => n10480, B1 => n9490, B2 => 
                           n10352, ZN => n1008);
   U1160 : OAI221_X1 port map( B1 => n8538, B2 => n9501, C1 => n8506, C2 => 
                           n9498, A => n954, ZN => n949);
   U1161 : AOI22_X1 port map( A1 => n9495, A2 => n10477, B1 => n9490, B2 => 
                           n10349, ZN => n954);
   U1162 : OAI221_X1 port map( B1 => n8855, B2 => n9453, C1 => n8823, C2 => 
                           n9450, A => n1016, ZN => n1011);
   U1163 : AOI22_X1 port map( A1 => n9447, A2 => n10576, B1 => n9442, B2 => 
                           n10016, ZN => n1016);
   U1164 : OAI221_X1 port map( B1 => n8516, B2 => n9499, C1 => n8484, C2 => 
                           n9496, A => n1350, ZN => n1345);
   U1165 : AOI22_X1 port map( A1 => n9493, A2 => n10499, B1 => n9492, B2 => 
                           n10371, ZN => n1350);
   U1166 : OAI221_X1 port map( B1 => n8832, B2 => n9451, C1 => n8800, C2 => 
                           n9448, A => n1430, ZN => n1425);
   U1167 : AOI22_X1 port map( A1 => n9445, A2 => n10007, B1 => n9444, B2 => 
                           n10039, ZN => n1430);
   U1168 : OAI221_X1 port map( B1 => n8534, B2 => n9501, C1 => n8502, C2 => 
                           n9498, A => n1026, ZN => n1021);
   U1169 : AOI22_X1 port map( A1 => n9495, A2 => n10481, B1 => n9490, B2 => 
                           n10353, ZN => n1026);
   U1170 : OAI221_X1 port map( B1 => n8539, B2 => n9501, C1 => n8507, C2 => 
                           n9498, A => n936, ZN => n931);
   U1171 : AOI22_X1 port map( A1 => n9495, A2 => n10476, B1 => n9490, B2 => 
                           n10348, ZN => n936);
   U1172 : OAI221_X1 port map( B1 => n8517, B2 => n9499, C1 => n8485, C2 => 
                           n9496, A => n1332, ZN => n1327);
   U1173 : AOI22_X1 port map( A1 => n9493, A2 => n10498, B1 => n9492, B2 => 
                           n10370, ZN => n1332);
   U1174 : OAI221_X1 port map( B1 => n8837, B2 => n9451, C1 => n8805, C2 => 
                           n9448, A => n1340, ZN => n1335);
   U1175 : AOI22_X1 port map( A1 => n9445, A2 => n10002, B1 => n9444, B2 => 
                           n10034, ZN => n1340);
   U1176 : OAI221_X1 port map( B1 => n8536, B2 => n9501, C1 => n8504, C2 => 
                           n9498, A => n990, ZN => n985);
   U1177 : AOI22_X1 port map( A1 => n9495, A2 => n10479, B1 => n9490, B2 => 
                           n10351, ZN => n990);
   U1178 : OAI221_X1 port map( B1 => n8856, B2 => n9453, C1 => n8824, C2 => 
                           n9450, A => n998, ZN => n993);
   U1179 : AOI22_X1 port map( A1 => n9447, A2 => n10575, B1 => n9442, B2 => 
                           n10015, ZN => n998);
   U1180 : OAI221_X1 port map( B1 => n8540, B2 => n9501, C1 => n8508, C2 => 
                           n9498, A => n918, ZN => n913);
   U1181 : AOI22_X1 port map( A1 => n9495, A2 => n10475, B1 => n9490, B2 => 
                           n10347, ZN => n918);
   U1182 : OAI221_X1 port map( B1 => n8518, B2 => n9499, C1 => n8486, C2 => 
                           n9496, A => n1314, ZN => n1309);
   U1183 : AOI22_X1 port map( A1 => n9493, A2 => n10497, B1 => n9491, B2 => 
                           n10369, ZN => n1314);
   U1184 : OAI221_X1 port map( B1 => n8838, B2 => n9451, C1 => n8806, C2 => 
                           n9448, A => n1322, ZN => n1317);
   U1185 : AOI22_X1 port map( A1 => n9445, A2 => n10001, B1 => n9443, B2 => 
                           n10033, ZN => n1322);
   U1186 : OAI221_X1 port map( B1 => n8860, B2 => n9453, C1 => n8828, C2 => 
                           n9450, A => n926, ZN => n921);
   U1187 : AOI22_X1 port map( A1 => n9447, A2 => n10571, B1 => n9442, B2 => 
                           n10011, ZN => n926);
   U1188 : OAI221_X1 port map( B1 => n8537, B2 => n9501, C1 => n8505, C2 => 
                           n9498, A => n972, ZN => n967);
   U1189 : AOI22_X1 port map( A1 => n9495, A2 => n10478, B1 => n9490, B2 => 
                           n10350, ZN => n972);
   U1190 : OAI221_X1 port map( B1 => n8519, B2 => n9499, C1 => n8487, C2 => 
                           n9496, A => n1296, ZN => n1291);
   U1191 : AOI22_X1 port map( A1 => n9493, A2 => n10496, B1 => n9491, B2 => 
                           n10368, ZN => n1296);
   U1192 : OAI221_X1 port map( B1 => n8857, B2 => n9453, C1 => n8825, C2 => 
                           n9450, A => n980, ZN => n975);
   U1193 : AOI22_X1 port map( A1 => n9447, A2 => n10574, B1 => n9442, B2 => 
                           n10014, ZN => n980);
   U1194 : OAI221_X1 port map( B1 => n8839, B2 => n9451, C1 => n8807, C2 => 
                           n9448, A => n1304, ZN => n1299);
   U1195 : AOI22_X1 port map( A1 => n9445, A2 => n10000, B1 => n9443, B2 => 
                           n10032, ZN => n1304);
   U1196 : OAI221_X1 port map( B1 => n8806, B2 => n9355, C1 => n8782, C2 => 
                           n9352, A => n1942, ZN => n1937);
   U1197 : AOI22_X1 port map( A1 => n9349, A2 => n10033, B1 => n9347, B2 => 
                           n10065, ZN => n1942);
   U1198 : OAI221_X1 port map( B1 => n8807, B2 => n9355, C1 => n8783, C2 => 
                           n9352, A => n1924, ZN => n1919);
   U1199 : AOI22_X1 port map( A1 => n9349, A2 => n10032, B1 => n9347, B2 => 
                           n10064, ZN => n1924);
   U1200 : OAI221_X1 port map( B1 => n8808, B2 => n9355, C1 => n8784, C2 => 
                           n9352, A => n1906, ZN => n1901);
   U1201 : AOI22_X1 port map( A1 => n9349, A2 => n10031, B1 => n9347, B2 => 
                           n10063, ZN => n1906);
   U1202 : OAI221_X1 port map( B1 => n8809, B2 => n9355, C1 => n8785, C2 => 
                           n9352, A => n1888, ZN => n1883);
   U1203 : AOI22_X1 port map( A1 => n9349, A2 => n10030, B1 => n9347, B2 => 
                           n10062, ZN => n1888);
   U1204 : OAI221_X1 port map( B1 => n8810, B2 => n9356, C1 => n8786, C2 => 
                           n9353, A => n1870, ZN => n1865);
   U1205 : AOI22_X1 port map( A1 => n9350, A2 => n10029, B1 => n9347, B2 => 
                           n10061, ZN => n1870);
   U1206 : OAI221_X1 port map( B1 => n8811, B2 => n9356, C1 => n8787, C2 => 
                           n9353, A => n1852, ZN => n1847);
   U1207 : AOI22_X1 port map( A1 => n9350, A2 => n10028, B1 => n9347, B2 => 
                           n10060, ZN => n1852);
   U1208 : OAI221_X1 port map( B1 => n8812, B2 => n9356, C1 => n8788, C2 => 
                           n9353, A => n1834, ZN => n1829);
   U1209 : AOI22_X1 port map( A1 => n9350, A2 => n10027, B1 => n9347, B2 => 
                           n10059, ZN => n1834);
   U1210 : OAI221_X1 port map( B1 => n8813, B2 => n9356, C1 => n8789, C2 => 
                           n9353, A => n1816, ZN => n1811);
   U1211 : AOI22_X1 port map( A1 => n9350, A2 => n10026, B1 => n9347, B2 => 
                           n10058, ZN => n1816);
   U1212 : OAI221_X1 port map( B1 => n8814, B2 => n9356, C1 => n8790, C2 => 
                           n9353, A => n1798, ZN => n1793);
   U1213 : AOI22_X1 port map( A1 => n9350, A2 => n10025, B1 => n9347, B2 => 
                           n10057, ZN => n1798);
   U1214 : OAI221_X1 port map( B1 => n8815, B2 => n9356, C1 => n8791, C2 => 
                           n9353, A => n1780, ZN => n1775);
   U1215 : AOI22_X1 port map( A1 => n9350, A2 => n10024, B1 => n9347, B2 => 
                           n10056, ZN => n1780);
   U1216 : OAI221_X1 port map( B1 => n8816, B2 => n9356, C1 => n8792, C2 => 
                           n9353, A => n1762, ZN => n1757);
   U1217 : AOI22_X1 port map( A1 => n9350, A2 => n10023, B1 => n9347, B2 => 
                           n10055, ZN => n1762);
   U1218 : OAI221_X1 port map( B1 => n8817, B2 => n9356, C1 => n8793, C2 => 
                           n9353, A => n1744, ZN => n1739);
   U1219 : AOI22_X1 port map( A1 => n9350, A2 => n10022, B1 => n9347, B2 => 
                           n10054, ZN => n1744);
   U1220 : OAI221_X1 port map( B1 => n8818, B2 => n9356, C1 => n8794, C2 => 
                           n9353, A => n1726, ZN => n1721);
   U1221 : AOI22_X1 port map( A1 => n9350, A2 => n10021, B1 => n9346, B2 => 
                           n10053, ZN => n1726);
   U1222 : OAI221_X1 port map( B1 => n8819, B2 => n9356, C1 => n8795, C2 => 
                           n9353, A => n1708, ZN => n1703);
   U1223 : AOI22_X1 port map( A1 => n9350, A2 => n10020, B1 => n9346, B2 => 
                           n10052, ZN => n1708);
   U1224 : OAI221_X1 port map( B1 => n8820, B2 => n9356, C1 => n8796, C2 => 
                           n9353, A => n1690, ZN => n1685);
   U1225 : AOI22_X1 port map( A1 => n9350, A2 => n10019, B1 => n9346, B2 => 
                           n10051, ZN => n1690);
   U1226 : OAI221_X1 port map( B1 => n8821, B2 => n9356, C1 => n8797, C2 => 
                           n9353, A => n1672, ZN => n1667);
   U1227 : AOI22_X1 port map( A1 => n9350, A2 => n10018, B1 => n9346, B2 => 
                           n10050, ZN => n1672);
   U1228 : OAI221_X1 port map( B1 => n8822, B2 => n9357, C1 => n8311, C2 => 
                           n9354, A => n1654, ZN => n1649);
   U1229 : AOI22_X1 port map( A1 => n9351, A2 => n10017, B1 => n9346, B2 => 
                           n10049, ZN => n1654);
   U1230 : OAI221_X1 port map( B1 => n8823, B2 => n9357, C1 => n8312, C2 => 
                           n9354, A => n1636, ZN => n1631);
   U1231 : AOI22_X1 port map( A1 => n9351, A2 => n10016, B1 => n9346, B2 => 
                           n10048, ZN => n1636);
   U1232 : OAI221_X1 port map( B1 => n8824, B2 => n9357, C1 => n8313, C2 => 
                           n9354, A => n1618, ZN => n1613);
   U1233 : AOI22_X1 port map( A1 => n9351, A2 => n10015, B1 => n9346, B2 => 
                           n10047, ZN => n1618);
   U1234 : OAI221_X1 port map( B1 => n8825, B2 => n9357, C1 => n8314, C2 => 
                           n9354, A => n1600, ZN => n1595);
   U1235 : AOI22_X1 port map( A1 => n9351, A2 => n10014, B1 => n9346, B2 => 
                           n10046, ZN => n1600);
   U1236 : OAI221_X1 port map( B1 => n8826, B2 => n9357, C1 => n8315, C2 => 
                           n9354, A => n1582, ZN => n1577);
   U1237 : AOI22_X1 port map( A1 => n9351, A2 => n10013, B1 => n9346, B2 => 
                           n10045, ZN => n1582);
   U1238 : OAI221_X1 port map( B1 => n8827, B2 => n9357, C1 => n8316, C2 => 
                           n9354, A => n1564, ZN => n1559);
   U1239 : AOI22_X1 port map( A1 => n9351, A2 => n10012, B1 => n9346, B2 => 
                           n10044, ZN => n1564);
   U1240 : OAI221_X1 port map( B1 => n8828, B2 => n9357, C1 => n8317, C2 => 
                           n9354, A => n1546, ZN => n1541);
   U1241 : AOI22_X1 port map( A1 => n9351, A2 => n10011, B1 => n9346, B2 => 
                           n10043, ZN => n1546);
   U1242 : OAI221_X1 port map( B1 => n8829, B2 => n9357, C1 => n8318, C2 => 
                           n9354, A => n1522, ZN => n1507);
   U1243 : AOI22_X1 port map( A1 => n9351, A2 => n10010, B1 => n9346, B2 => 
                           n10042, ZN => n1522);
   U1244 : OAI221_X1 port map( B1 => n8922, B2 => n9439, C1 => n8890, C2 => 
                           n9436, A => n1395, ZN => n1388);
   U1245 : AOI22_X1 port map( A1 => n9433, A2 => n10341, B1 => n9432, B2 => 
                           n9949, ZN => n1395);
   U1246 : OAI221_X1 port map( B1 => n8923, B2 => n9439, C1 => n8891, C2 => 
                           n9436, A => n1377, ZN => n1370);
   U1247 : AOI22_X1 port map( A1 => n9433, A2 => n10340, B1 => n9432, B2 => 
                           n9948, ZN => n1377);
   U1248 : OAI221_X1 port map( B1 => n2247, B2 => n9488, C1 => n8388, C2 => 
                           n9485, A => n1225, ZN => n1218);
   U1249 : AOI22_X1 port map( A1 => n9482, A2 => n10212, B1 => n9479, B2 => 
                           n10644, ZN => n1225);
   U1250 : OAI221_X1 port map( B1 => n2239, B2 => n9488, C1 => n8389, C2 => 
                           n9485, A => n1207, ZN => n1200);
   U1251 : AOI22_X1 port map( A1 => n9482, A2 => n10211, B1 => n9479, B2 => 
                           n10643, ZN => n1207);
   U1252 : OAI221_X1 port map( B1 => n2231, B2 => n9488, C1 => n8390, C2 => 
                           n9485, A => n1189, ZN => n1182);
   U1253 : AOI22_X1 port map( A1 => n9482, A2 => n10210, B1 => n9479, B2 => 
                           n10642, ZN => n1189);
   U1254 : OAI221_X1 port map( B1 => n2191, B2 => n9488, C1 => n8395, C2 => 
                           n9485, A => n1099, ZN => n1092);
   U1255 : AOI22_X1 port map( A1 => n9482, A2 => n10205, B1 => n9478, B2 => 
                           n10637, ZN => n1099);
   U1256 : OAI221_X1 port map( B1 => n2271, B2 => n9487, C1 => n8385, C2 => 
                           n9484, A => n1279, ZN => n1272);
   U1257 : AOI22_X1 port map( A1 => n9481, A2 => n10215, B1 => n9479, B2 => 
                           n10647, ZN => n1279);
   U1258 : OAI221_X1 port map( B1 => n2263, B2 => n9487, C1 => n8386, C2 => 
                           n9484, A => n1261, ZN => n1254);
   U1259 : AOI22_X1 port map( A1 => n9481, A2 => n10214, B1 => n9479, B2 => 
                           n10646, ZN => n1261);
   U1260 : OAI221_X1 port map( B1 => n2175, B2 => n9488, C1 => n8397, C2 => 
                           n9485, A => n1063, ZN => n1056);
   U1261 : AOI22_X1 port map( A1 => n9482, A2 => n10203, B1 => n9478, B2 => 
                           n10635, ZN => n1063);
   U1262 : OAI221_X1 port map( B1 => n2183, B2 => n9488, C1 => n8396, C2 => 
                           n9485, A => n1081, ZN => n1074);
   U1263 : AOI22_X1 port map( A1 => n9482, A2 => n10204, B1 => n9478, B2 => 
                           n10636, ZN => n1081);
   U1264 : OAI221_X1 port map( B1 => n8938, B2 => n9440, C1 => n8906, C2 => 
                           n9437, A => n1107, ZN => n1100);
   U1265 : AOI22_X1 port map( A1 => n9434, A2 => n10325, B1 => n9430, B2 => 
                           n9933, ZN => n1107);
   U1266 : OAI221_X1 port map( B1 => n8933, B2 => n9440, C1 => n8901, C2 => 
                           n9437, A => n1197, ZN => n1190);
   U1267 : AOI22_X1 port map( A1 => n9434, A2 => n10330, B1 => n9431, B2 => 
                           n9938, ZN => n1197);
   U1268 : OAI221_X1 port map( B1 => n8939, B2 => n9440, C1 => n8907, C2 => 
                           n9437, A => n1089, ZN => n1082);
   U1269 : AOI22_X1 port map( A1 => n9434, A2 => n10324, B1 => n9430, B2 => 
                           n9932, ZN => n1089);
   U1270 : OAI221_X1 port map( B1 => n8929, B2 => n9439, C1 => n8897, C2 => 
                           n9436, A => n1269, ZN => n1262);
   U1271 : AOI22_X1 port map( A1 => n9433, A2 => n10334, B1 => n9431, B2 => 
                           n9942, ZN => n1269);
   U1272 : OAI221_X1 port map( B1 => n8940, B2 => n9440, C1 => n8908, C2 => 
                           n9437, A => n1071, ZN => n1064);
   U1273 : AOI22_X1 port map( A1 => n9434, A2 => n10323, B1 => n9430, B2 => 
                           n9931, ZN => n1071);
   U1274 : OAI221_X1 port map( B1 => n2223, B2 => n9488, C1 => n8391, C2 => 
                           n9485, A => n1171, ZN => n1164);
   U1275 : AOI22_X1 port map( A1 => n9482, A2 => n10209, B1 => n9479, B2 => 
                           n10641, ZN => n1171);
   U1276 : OAI221_X1 port map( B1 => n2255, B2 => n9488, C1 => n8387, C2 => 
                           n9485, A => n1243, ZN => n1236);
   U1277 : AOI22_X1 port map( A1 => n9482, A2 => n10213, B1 => n9479, B2 => 
                           n10645, ZN => n1243);
   U1278 : OAI221_X1 port map( B1 => n2167, B2 => n9488, C1 => n8398, C2 => 
                           n9485, A => n1045, ZN => n1038);
   U1279 : AOI22_X1 port map( A1 => n9482, A2 => n10202, B1 => n9478, B2 => 
                           n10634, ZN => n1045);
   U1280 : OAI221_X1 port map( B1 => n8934, B2 => n9440, C1 => n8902, C2 => 
                           n9437, A => n1179, ZN => n1172);
   U1281 : AOI22_X1 port map( A1 => n9434, A2 => n10329, B1 => n9431, B2 => 
                           n9937, ZN => n1179);
   U1282 : OAI221_X1 port map( B1 => n8930, B2 => n9440, C1 => n8898, C2 => 
                           n9437, A => n1251, ZN => n1244);
   U1283 : AOI22_X1 port map( A1 => n9434, A2 => n10333, B1 => n9431, B2 => 
                           n9941, ZN => n1251);
   U1284 : OAI221_X1 port map( B1 => n8941, B2 => n9440, C1 => n8909, C2 => 
                           n9437, A => n1053, ZN => n1046);
   U1285 : AOI22_X1 port map( A1 => n9434, A2 => n10322, B1 => n9430, B2 => 
                           n9930, ZN => n1053);
   U1286 : OAI221_X1 port map( B1 => n2215, B2 => n9488, C1 => n8392, C2 => 
                           n9485, A => n1153, ZN => n1146);
   U1287 : AOI22_X1 port map( A1 => n9482, A2 => n10208, B1 => n9479, B2 => 
                           n10640, ZN => n1153);
   U1288 : OAI221_X1 port map( B1 => n2207, B2 => n9488, C1 => n8393, C2 => 
                           n9485, A => n1135, ZN => n1128);
   U1289 : AOI22_X1 port map( A1 => n9482, A2 => n10207, B1 => n9479, B2 => 
                           n10639, ZN => n1135);
   U1290 : OAI221_X1 port map( B1 => n2199, B2 => n9488, C1 => n8394, C2 => 
                           n9485, A => n1117, ZN => n1110);
   U1291 : AOI22_X1 port map( A1 => n9482, A2 => n10206, B1 => n9479, B2 => 
                           n10638, ZN => n1117);
   U1292 : OAI221_X1 port map( B1 => n8937, B2 => n9440, C1 => n8905, C2 => 
                           n9437, A => n1125, ZN => n1118);
   U1293 : AOI22_X1 port map( A1 => n9434, A2 => n10326, B1 => n9431, B2 => 
                           n9934, ZN => n1125);
   U1294 : OAI221_X1 port map( B1 => n8919, B2 => n9439, C1 => n8887, C2 => 
                           n9436, A => n1449, ZN => n1442);
   U1295 : AOI22_X1 port map( A1 => n9433, A2 => n10344, B1 => n9432, B2 => 
                           n9952, ZN => n1449);
   U1296 : OAI221_X1 port map( B1 => n8920, B2 => n9439, C1 => n8888, C2 => 
                           n9436, A => n1431, ZN => n1424);
   U1297 : AOI22_X1 port map( A1 => n9433, A2 => n10343, B1 => n9432, B2 => 
                           n9951, ZN => n1431);
   U1298 : OAI221_X1 port map( B1 => n8943, B2 => n9441, C1 => n8911, C2 => 
                           n9438, A => n1017, ZN => n1010);
   U1299 : AOI22_X1 port map( A1 => n9435, A2 => n10568, B1 => n9430, B2 => 
                           n9928, ZN => n1017);
   U1300 : OAI221_X1 port map( B1 => n8925, B2 => n9439, C1 => n8893, C2 => 
                           n9436, A => n1341, ZN => n1334);
   U1301 : AOI22_X1 port map( A1 => n9433, A2 => n10338, B1 => n9432, B2 => 
                           n9946, ZN => n1341);
   U1302 : OAI221_X1 port map( B1 => n2287, B2 => n9487, C1 => n8383, C2 => 
                           n9484, A => n1315, ZN => n1308);
   U1303 : AOI22_X1 port map( A1 => n9481, A2 => n10217, B1 => n9479, B2 => 
                           n10649, ZN => n1315);
   U1304 : OAI221_X1 port map( B1 => n8944, B2 => n9441, C1 => n8912, C2 => 
                           n9438, A => n999, ZN => n992);
   U1305 : AOI22_X1 port map( A1 => n9435, A2 => n10567, B1 => n9430, B2 => 
                           n9927, ZN => n999);
   U1306 : OAI221_X1 port map( B1 => n2279, B2 => n9487, C1 => n8384, C2 => 
                           n9484, A => n1297, ZN => n1290);
   U1307 : AOI22_X1 port map( A1 => n9481, A2 => n10216, B1 => n9479, B2 => 
                           n10648, ZN => n1297);
   U1308 : OAI221_X1 port map( B1 => n8926, B2 => n9439, C1 => n8894, C2 => 
                           n9436, A => n1323, ZN => n1316);
   U1309 : AOI22_X1 port map( A1 => n9433, A2 => n10337, B1 => n9431, B2 => 
                           n9945, ZN => n1323);
   U1310 : OAI221_X1 port map( B1 => n8948, B2 => n9441, C1 => n8916, C2 => 
                           n9438, A => n927, ZN => n920);
   U1311 : AOI22_X1 port map( A1 => n9435, A2 => n10563, B1 => n9430, B2 => 
                           n9923, ZN => n927);
   U1312 : OAI221_X1 port map( B1 => n8945, B2 => n9441, C1 => n8913, C2 => 
                           n9438, A => n981, ZN => n974);
   U1313 : AOI22_X1 port map( A1 => n9435, A2 => n10566, B1 => n9430, B2 => 
                           n9926, ZN => n981);
   U1314 : OAI221_X1 port map( B1 => n8927, B2 => n9439, C1 => n8895, C2 => 
                           n9436, A => n1305, ZN => n1298);
   U1315 : AOI22_X1 port map( A1 => n9433, A2 => n10336, B1 => n9431, B2 => 
                           n9944, ZN => n1305);
   U1316 : OAI221_X1 port map( B1 => n8894, B2 => n9343, C1 => n8870, C2 => 
                           n9340, A => n1943, ZN => n1936);
   U1317 : AOI22_X1 port map( A1 => n9337, A2 => n9945, B1 => n9335, B2 => 
                           n9977, ZN => n1943);
   U1318 : OAI221_X1 port map( B1 => n8895, B2 => n9343, C1 => n8871, C2 => 
                           n9340, A => n1925, ZN => n1918);
   U1319 : AOI22_X1 port map( A1 => n9337, A2 => n9944, B1 => n9335, B2 => 
                           n9976, ZN => n1925);
   U1320 : OAI221_X1 port map( B1 => n8896, B2 => n9343, C1 => n8872, C2 => 
                           n9340, A => n1907, ZN => n1900);
   U1321 : AOI22_X1 port map( A1 => n9337, A2 => n9943, B1 => n9335, B2 => 
                           n9975, ZN => n1907);
   U1322 : OAI221_X1 port map( B1 => n8897, B2 => n9343, C1 => n8873, C2 => 
                           n9340, A => n1889, ZN => n1882);
   U1323 : AOI22_X1 port map( A1 => n9337, A2 => n9942, B1 => n9335, B2 => 
                           n9974, ZN => n1889);
   U1324 : OAI221_X1 port map( B1 => n8898, B2 => n9344, C1 => n8874, C2 => 
                           n9341, A => n1871, ZN => n1864);
   U1325 : AOI22_X1 port map( A1 => n9338, A2 => n9941, B1 => n9335, B2 => 
                           n9973, ZN => n1871);
   U1326 : OAI221_X1 port map( B1 => n8899, B2 => n9344, C1 => n8875, C2 => 
                           n9341, A => n1853, ZN => n1846);
   U1327 : AOI22_X1 port map( A1 => n9338, A2 => n9940, B1 => n9335, B2 => 
                           n9972, ZN => n1853);
   U1328 : OAI221_X1 port map( B1 => n8900, B2 => n9344, C1 => n8876, C2 => 
                           n9341, A => n1835, ZN => n1828);
   U1329 : AOI22_X1 port map( A1 => n9338, A2 => n9939, B1 => n9335, B2 => 
                           n9971, ZN => n1835);
   U1330 : OAI221_X1 port map( B1 => n8901, B2 => n9344, C1 => n8877, C2 => 
                           n9341, A => n1817, ZN => n1810);
   U1331 : AOI22_X1 port map( A1 => n9338, A2 => n9938, B1 => n9335, B2 => 
                           n9970, ZN => n1817);
   U1332 : OAI221_X1 port map( B1 => n8902, B2 => n9344, C1 => n8878, C2 => 
                           n9341, A => n1799, ZN => n1792);
   U1333 : AOI22_X1 port map( A1 => n9338, A2 => n9937, B1 => n9335, B2 => 
                           n9969, ZN => n1799);
   U1334 : OAI221_X1 port map( B1 => n8903, B2 => n9344, C1 => n8879, C2 => 
                           n9341, A => n1781, ZN => n1774);
   U1335 : AOI22_X1 port map( A1 => n9338, A2 => n9936, B1 => n9335, B2 => 
                           n9968, ZN => n1781);
   U1336 : OAI221_X1 port map( B1 => n8904, B2 => n9344, C1 => n8880, C2 => 
                           n9341, A => n1763, ZN => n1756);
   U1337 : AOI22_X1 port map( A1 => n9338, A2 => n9935, B1 => n9335, B2 => 
                           n9967, ZN => n1763);
   U1338 : OAI221_X1 port map( B1 => n8905, B2 => n9344, C1 => n8881, C2 => 
                           n9341, A => n1745, ZN => n1738);
   U1339 : AOI22_X1 port map( A1 => n9338, A2 => n9934, B1 => n9335, B2 => 
                           n9966, ZN => n1745);
   U1340 : OAI221_X1 port map( B1 => n8906, B2 => n9344, C1 => n8882, C2 => 
                           n9341, A => n1727, ZN => n1720);
   U1341 : AOI22_X1 port map( A1 => n9338, A2 => n9933, B1 => n9334, B2 => 
                           n9965, ZN => n1727);
   U1342 : OAI221_X1 port map( B1 => n8907, B2 => n9344, C1 => n8883, C2 => 
                           n9341, A => n1709, ZN => n1702);
   U1343 : AOI22_X1 port map( A1 => n9338, A2 => n9932, B1 => n9334, B2 => 
                           n9964, ZN => n1709);
   U1344 : OAI221_X1 port map( B1 => n8908, B2 => n9344, C1 => n8884, C2 => 
                           n9341, A => n1691, ZN => n1684);
   U1345 : AOI22_X1 port map( A1 => n9338, A2 => n9931, B1 => n9334, B2 => 
                           n9963, ZN => n1691);
   U1346 : OAI221_X1 port map( B1 => n8909, B2 => n9344, C1 => n8885, C2 => 
                           n9341, A => n1673, ZN => n1666);
   U1347 : AOI22_X1 port map( A1 => n9338, A2 => n9930, B1 => n9334, B2 => 
                           n9962, ZN => n1673);
   U1348 : OAI221_X1 port map( B1 => n8910, B2 => n9345, C1 => n8303, C2 => 
                           n9342, A => n1655, ZN => n1648);
   U1349 : AOI22_X1 port map( A1 => n9339, A2 => n9929, B1 => n9334, B2 => 
                           n9961, ZN => n1655);
   U1350 : OAI221_X1 port map( B1 => n8911, B2 => n9345, C1 => n8304, C2 => 
                           n9342, A => n1637, ZN => n1630);
   U1351 : AOI22_X1 port map( A1 => n9339, A2 => n9928, B1 => n9334, B2 => 
                           n9960, ZN => n1637);
   U1352 : OAI221_X1 port map( B1 => n8912, B2 => n9345, C1 => n8305, C2 => 
                           n9342, A => n1619, ZN => n1612);
   U1353 : AOI22_X1 port map( A1 => n9339, A2 => n9927, B1 => n9334, B2 => 
                           n9959, ZN => n1619);
   U1354 : OAI221_X1 port map( B1 => n8913, B2 => n9345, C1 => n8306, C2 => 
                           n9342, A => n1601, ZN => n1594);
   U1355 : AOI22_X1 port map( A1 => n9339, A2 => n9926, B1 => n9334, B2 => 
                           n9958, ZN => n1601);
   U1356 : OAI221_X1 port map( B1 => n8914, B2 => n9345, C1 => n8307, C2 => 
                           n9342, A => n1583, ZN => n1576);
   U1357 : AOI22_X1 port map( A1 => n9339, A2 => n9925, B1 => n9334, B2 => 
                           n9957, ZN => n1583);
   U1358 : OAI221_X1 port map( B1 => n8915, B2 => n9345, C1 => n8308, C2 => 
                           n9342, A => n1565, ZN => n1558);
   U1359 : AOI22_X1 port map( A1 => n9339, A2 => n9924, B1 => n9334, B2 => 
                           n9956, ZN => n1565);
   U1360 : OAI221_X1 port map( B1 => n8916, B2 => n9345, C1 => n8309, C2 => 
                           n9342, A => n1547, ZN => n1540);
   U1361 : AOI22_X1 port map( A1 => n9339, A2 => n9923, B1 => n9334, B2 => 
                           n9955, ZN => n1547);
   U1362 : OAI221_X1 port map( B1 => n8917, B2 => n9345, C1 => n8310, C2 => 
                           n9342, A => n1527, ZN => n1506);
   U1363 : AOI22_X1 port map( A1 => n9339, A2 => n9922, B1 => n9334, B2 => 
                           n9954, ZN => n1527);
   U1364 : AOI22_X1 port map( A1 => n9458, A2 => n10124, B1 => n9455, B2 => 
                           n10156, ZN => n1231);
   U1365 : AOI22_X1 port map( A1 => n9457, A2 => n10137, B1 => n9456, B2 => 
                           n10169, ZN => n1476);
   U1366 : AOI22_X1 port map( A1 => n9458, A2 => n10120, B1 => n9455, B2 => 
                           n10152, ZN => n1159);
   U1367 : AOI22_X1 port map( A1 => n9457, A2 => n10131, B1 => n9456, B2 => 
                           n10163, ZN => n1357);
   U1368 : AOI22_X1 port map( A1 => n9470, A2 => n10180, B1 => n9467, B2 => 
                           n10244, ZN => n1230);
   U1369 : AOI22_X1 port map( A1 => n9469, A2 => n10193, B1 => n9468, B2 => 
                           n10257, ZN => n1475);
   U1370 : AOI22_X1 port map( A1 => n9470, A2 => n10176, B1 => n9467, B2 => 
                           n10240, ZN => n1158);
   U1371 : AOI22_X1 port map( A1 => n9469, A2 => n10187, B1 => n9468, B2 => 
                           n10251, ZN => n1356);
   U1372 : NOR4_X1 port map( A1 => n1452, A2 => n1453, A3 => n1454, A4 => n1455
                           , ZN => n1451);
   U1373 : OAI221_X1 port map( B1 => n8918, B2 => n9439, C1 => n8886, C2 => 
                           n9436, A => n1479, ZN => n1471);
   U1374 : NOR4_X1 port map( A1 => n1218, A2 => n1219, A3 => n1220, A4 => n1221
                           , ZN => n1217);
   U1375 : OAI221_X1 port map( B1 => n8931, B2 => n9440, C1 => n8899, C2 => 
                           n9437, A => n1233, ZN => n1226);
   U1376 : NOR4_X1 port map( A1 => n1146, A2 => n1147, A3 => n1148, A4 => n1149
                           , ZN => n1145);
   U1377 : OAI221_X1 port map( B1 => n8935, B2 => n9440, C1 => n8903, C2 => 
                           n9437, A => n1161, ZN => n1154);
   U1378 : NOR4_X1 port map( A1 => n1308, A2 => n1309, A3 => n1310, A4 => n1311
                           , ZN => n1307);
   U1379 : NOR4_X1 port map( A1 => n1316, A2 => n1317, A3 => n1318, A4 => n1319
                           , ZN => n1306);
   U1380 : OAI221_X1 port map( B1 => n8247, B2 => n9511, C1 => n8228, C2 => 
                           n9508, A => n1313, ZN => n1310);
   U1381 : OAI221_X1 port map( B1 => n8921, B2 => n9439, C1 => n8889, C2 => 
                           n9436, A => n1413, ZN => n1406);
   U1382 : AOI22_X1 port map( A1 => n9433, A2 => n10342, B1 => n9432, B2 => 
                           n9950, ZN => n1413);
   U1383 : OAI221_X1 port map( B1 => n8949, B2 => n9441, C1 => n8917, C2 => 
                           n9438, A => n907, ZN => n886);
   U1384 : AOI22_X1 port map( A1 => n9435, A2 => n10562, B1 => n9430, B2 => 
                           n9922, ZN => n907);
   U1385 : OAI221_X1 port map( B1 => n8932, B2 => n9440, C1 => n8900, C2 => 
                           n9437, A => n1215, ZN => n1208);
   U1386 : AOI22_X1 port map( A1 => n9434, A2 => n10331, B1 => n9431, B2 => 
                           n9939, ZN => n1215);
   U1387 : OAI221_X1 port map( B1 => n8928, B2 => n9439, C1 => n8896, C2 => 
                           n9436, A => n1287, ZN => n1280);
   U1388 : AOI22_X1 port map( A1 => n9433, A2 => n10335, B1 => n9431, B2 => 
                           n9943, ZN => n1287);
   U1389 : OAI221_X1 port map( B1 => n8936, B2 => n9440, C1 => n8904, C2 => 
                           n9437, A => n1143, ZN => n1136);
   U1390 : AOI22_X1 port map( A1 => n9434, A2 => n10327, B1 => n9431, B2 => 
                           n9935, ZN => n1143);
   U1391 : OAI221_X1 port map( B1 => n8946, B2 => n9441, C1 => n8914, C2 => 
                           n9438, A => n963, ZN => n956);
   U1392 : AOI22_X1 port map( A1 => n9435, A2 => n10565, B1 => n9430, B2 => 
                           n9925, ZN => n963);
   U1393 : OAI221_X1 port map( B1 => n8942, B2 => n9441, C1 => n8910, C2 => 
                           n9438, A => n1035, ZN => n1028);
   U1394 : AOI22_X1 port map( A1 => n9435, A2 => n10569, B1 => n9430, B2 => 
                           n9929, ZN => n1035);
   U1395 : OAI221_X1 port map( B1 => n8947, B2 => n9441, C1 => n8915, C2 => 
                           n9438, A => n945, ZN => n938);
   U1396 : AOI22_X1 port map( A1 => n9435, A2 => n10564, B1 => n9430, B2 => 
                           n9924, ZN => n945);
   U1397 : AND3_X1 port map( A1 => ADD_RD2(4), A2 => n10662, A3 => RD2, ZN => 
                           n2088);
   U1398 : OAI221_X1 port map( B1 => n8833, B2 => n9451, C1 => n8801, C2 => 
                           n9448, A => n1412, ZN => n1407);
   U1399 : AOI22_X1 port map( A1 => n9445, A2 => n10006, B1 => n9444, B2 => 
                           n10038, ZN => n1412);
   U1400 : OAI221_X1 port map( B1 => n8861, B2 => n9453, C1 => n8829, C2 => 
                           n9450, A => n902, ZN => n887);
   U1401 : AOI22_X1 port map( A1 => n9447, A2 => n10570, B1 => n9442, B2 => 
                           n10010, ZN => n902);
   U1402 : OAI221_X1 port map( B1 => n8843, B2 => n9452, C1 => n8811, C2 => 
                           n9449, A => n1232, ZN => n1227);
   U1403 : AOI22_X1 port map( A1 => n9446, A2 => n9996, B1 => n9443, B2 => 
                           n10028, ZN => n1232);
   U1404 : OAI221_X1 port map( B1 => n8830, B2 => n9451, C1 => n8798, C2 => 
                           n9448, A => n1478, ZN => n1472);
   U1405 : AOI22_X1 port map( A1 => n9445, A2 => n10009, B1 => n9444, B2 => 
                           n10041, ZN => n1478);
   U1406 : OAI221_X1 port map( B1 => n8844, B2 => n9452, C1 => n8812, C2 => 
                           n9449, A => n1214, ZN => n1209);
   U1407 : AOI22_X1 port map( A1 => n9446, A2 => n9995, B1 => n9443, B2 => 
                           n10027, ZN => n1214);
   U1408 : OAI221_X1 port map( B1 => n8840, B2 => n9451, C1 => n8808, C2 => 
                           n9448, A => n1286, ZN => n1281);
   U1409 : AOI22_X1 port map( A1 => n9445, A2 => n9999, B1 => n9443, B2 => 
                           n10031, ZN => n1286);
   U1410 : OAI221_X1 port map( B1 => n8847, B2 => n9452, C1 => n8815, C2 => 
                           n9449, A => n1160, ZN => n1155);
   U1411 : AOI22_X1 port map( A1 => n9446, A2 => n9992, B1 => n9443, B2 => 
                           n10024, ZN => n1160);
   U1412 : OAI221_X1 port map( B1 => n8848, B2 => n9452, C1 => n8816, C2 => 
                           n9449, A => n1142, ZN => n1137);
   U1413 : AOI22_X1 port map( A1 => n9446, A2 => n9991, B1 => n9443, B2 => 
                           n10023, ZN => n1142);
   U1414 : OAI221_X1 port map( B1 => n8858, B2 => n9453, C1 => n8826, C2 => 
                           n9450, A => n962, ZN => n957);
   U1415 : AOI22_X1 port map( A1 => n9447, A2 => n10573, B1 => n9442, B2 => 
                           n10013, ZN => n962);
   U1416 : OAI221_X1 port map( B1 => n8836, B2 => n9451, C1 => n8804, C2 => 
                           n9448, A => n1358, ZN => n1353);
   U1417 : AOI22_X1 port map( A1 => n9445, A2 => n10003, B1 => n9444, B2 => 
                           n10035, ZN => n1358);
   U1418 : OAI221_X1 port map( B1 => n8854, B2 => n9453, C1 => n8822, C2 => 
                           n9450, A => n1034, ZN => n1029);
   U1419 : AOI22_X1 port map( A1 => n9447, A2 => n10577, B1 => n9442, B2 => 
                           n10017, ZN => n1034);
   U1420 : OAI221_X1 port map( B1 => n8859, B2 => n9453, C1 => n8827, C2 => 
                           n9450, A => n944, ZN => n939);
   U1421 : AOI22_X1 port map( A1 => n9447, A2 => n10572, B1 => n9442, B2 => 
                           n10012, ZN => n944);
   U1422 : OAI221_X1 port map( B1 => n8777, B2 => n9463, C1 => n8239, C2 => 
                           n9460, A => n1411, ZN => n1408);
   U1423 : AOI22_X1 port map( A1 => n9457, A2 => n10134, B1 => n9456, B2 => 
                           n10166, ZN => n1411);
   U1424 : OAI221_X1 port map( B1 => n8318, B2 => n9465, C1 => n8183, C2 => 
                           n9462, A => n897, ZN => n888);
   U1425 : AOI22_X1 port map( A1 => n9459, A2 => n10106, B1 => n9454, B2 => 
                           n10138, ZN => n897);
   U1426 : OAI221_X1 port map( B1 => n8788, B2 => n9464, C1 => n8217, C2 => 
                           n9461, A => n1213, ZN => n1210);
   U1427 : AOI22_X1 port map( A1 => n9458, A2 => n10123, B1 => n9455, B2 => 
                           n10155, ZN => n1213);
   U1428 : OAI221_X1 port map( B1 => n8784, B2 => n9463, C1 => n8225, C2 => 
                           n9460, A => n1285, ZN => n1282);
   U1429 : AOI22_X1 port map( A1 => n9457, A2 => n10127, B1 => n9455, B2 => 
                           n10159, ZN => n1285);
   U1430 : OAI221_X1 port map( B1 => n8792, B2 => n9464, C1 => n8209, C2 => 
                           n9461, A => n1141, ZN => n1138);
   U1431 : AOI22_X1 port map( A1 => n9458, A2 => n10119, B1 => n9455, B2 => 
                           n10151, ZN => n1141);
   U1432 : OAI221_X1 port map( B1 => n8315, B2 => n9465, C1 => n8189, C2 => 
                           n9462, A => n961, ZN => n958);
   U1433 : AOI22_X1 port map( A1 => n9459, A2 => n10109, B1 => n9454, B2 => 
                           n10141, ZN => n961);
   U1434 : OAI221_X1 port map( B1 => n8311, B2 => n9465, C1 => n8197, C2 => 
                           n9462, A => n1033, ZN => n1030);
   U1435 : AOI22_X1 port map( A1 => n9459, A2 => n10113, B1 => n9454, B2 => 
                           n10145, ZN => n1033);
   U1436 : OAI221_X1 port map( B1 => n8316, B2 => n9465, C1 => n8187, C2 => 
                           n9462, A => n943, ZN => n940);
   U1437 : AOI22_X1 port map( A1 => n9459, A2 => n10108, B1 => n9454, B2 => 
                           n10140, ZN => n943);
   U1438 : OAI221_X1 port map( B1 => n8657, B2 => n9475, C1 => n8633, C2 => 
                           n9472, A => n1410, ZN => n1409);
   U1439 : AOI22_X1 port map( A1 => n9469, A2 => n10190, B1 => n9468, B2 => 
                           n10254, ZN => n1410);
   U1440 : OAI221_X1 port map( B1 => n8685, B2 => n9477, C1 => n8302, C2 => 
                           n9474, A => n892, ZN => n889);
   U1441 : AOI22_X1 port map( A1 => n9471, A2 => n10578, B1 => n9466, B2 => 
                           n10226, ZN => n892);
   U1442 : OAI221_X1 port map( B1 => n8668, B2 => n9476, C1 => n8644, C2 => 
                           n9473, A => n1212, ZN => n1211);
   U1443 : AOI22_X1 port map( A1 => n9470, A2 => n10179, B1 => n9467, B2 => 
                           n10243, ZN => n1212);
   U1444 : OAI221_X1 port map( B1 => n8664, B2 => n9475, C1 => n8640, C2 => 
                           n9472, A => n1284, ZN => n1283);
   U1445 : AOI22_X1 port map( A1 => n9469, A2 => n10183, B1 => n9467, B2 => 
                           n10247, ZN => n1284);
   U1446 : OAI221_X1 port map( B1 => n8672, B2 => n9476, C1 => n8648, C2 => 
                           n9473, A => n1140, ZN => n1139);
   U1447 : AOI22_X1 port map( A1 => n9470, A2 => n10175, B1 => n9467, B2 => 
                           n10239, ZN => n1140);
   U1448 : OAI221_X1 port map( B1 => n8682, B2 => n9477, C1 => n8299, C2 => 
                           n9474, A => n960, ZN => n959);
   U1449 : AOI22_X1 port map( A1 => n9471, A2 => n10581, B1 => n9466, B2 => 
                           n10229, ZN => n960);
   U1450 : OAI221_X1 port map( B1 => n8678, B2 => n9477, C1 => n8295, C2 => 
                           n9474, A => n1032, ZN => n1031);
   U1451 : AOI22_X1 port map( A1 => n9471, A2 => n10585, B1 => n9466, B2 => 
                           n10233, ZN => n1032);
   U1452 : OAI221_X1 port map( B1 => n8683, B2 => n9477, C1 => n8300, C2 => 
                           n9474, A => n942, ZN => n941);
   U1453 : AOI22_X1 port map( A1 => n9471, A2 => n10580, B1 => n9466, B2 => 
                           n10228, ZN => n942);
   U1454 : AND3_X1 port map( A1 => RD2, A2 => ADD_RD2(4), A3 => ADD_RD2(3), ZN 
                           => n2077);
   U1455 : AND3_X1 port map( A1 => RD2, A2 => n10661, A3 => ADD_RD2(3), ZN => 
                           n2095);
   U1456 : AND3_X1 port map( A1 => n10662, A2 => n10661, A3 => RD2, ZN => n2098
                           );
   U1457 : OAI22_X1 port map( A1 => n9870, A2 => n9259, B1 => n2157, B2 => 
                           n9867, ZN => n9198);
   U1458 : OAI22_X1 port map( A1 => n9870, A2 => n9256, B1 => n2149, B2 => 
                           n9868, ZN => n9199);
   U1459 : OAI22_X1 port map( A1 => n9870, A2 => n9253, B1 => n2141, B2 => 
                           n9867, ZN => n9200);
   U1460 : OAI22_X1 port map( A1 => n9869, A2 => n9250, B1 => n2133, B2 => 
                           n9868, ZN => n9201);
   U1461 : OAI22_X1 port map( A1 => n9869, A2 => n9247, B1 => n2125, B2 => 
                           n9867, ZN => n9202);
   U1462 : OAI22_X1 port map( A1 => n9869, A2 => n9244, B1 => n2117, B2 => 
                           n9868, ZN => n9203);
   U1463 : OAI22_X1 port map( A1 => n9869, A2 => n9241, B1 => n2109, B2 => 
                           n9867, ZN => n9204);
   U1464 : OAI22_X1 port map( A1 => n9869, A2 => n9238, B1 => n2101, B2 => 
                           n9868, ZN => n9205);
   U1465 : OAI221_X1 port map( B1 => n2327, B2 => n9487, C1 => n8378, C2 => 
                           n9484, A => n1405, ZN => n1398);
   U1466 : AOI22_X1 port map( A1 => n9481, A2 => n10222, B1 => n9480, B2 => 
                           n10654, ZN => n1405);
   U1467 : AOI22_X1 port map( A1 => n9505, A2 => n10606, B1 => n9504, B2 => 
                           n10438, ZN => n1403);
   U1468 : OAI221_X1 port map( B1 => n8629, B2 => n9525, C1 => n8597, C2 => 
                           n9522, A => n868, ZN => n865);
   U1469 : AOI22_X1 port map( A1 => n9519, A2 => n10442, B1 => n9514, B2 => 
                           n10258, ZN => n868);
   U1470 : OAI221_X1 port map( B1 => n2319, B2 => n9487, C1 => n8379, C2 => 
                           n9484, A => n1387, ZN => n1380);
   U1471 : AOI22_X1 port map( A1 => n9481, A2 => n10221, B1 => n9480, B2 => 
                           n10653, ZN => n1387);
   U1472 : AOI22_X1 port map( A1 => n9505, A2 => n10605, B1 => n9504, B2 => 
                           n10437, ZN => n1385);
   U1473 : OAI221_X1 port map( B1 => n2311, B2 => n9487, C1 => n8380, C2 => 
                           n9484, A => n1369, ZN => n1362);
   U1474 : AOI22_X1 port map( A1 => n9481, A2 => n10220, B1 => n9480, B2 => 
                           n10652, ZN => n1369);
   U1475 : AOI22_X1 port map( A1 => n9505, A2 => n10604, B1 => n9504, B2 => 
                           n10436, ZN => n1367);
   U1476 : OAI221_X1 port map( B1 => n8611, B2 => n9524, C1 => n8579, C2 => 
                           n9521, A => n1222, ZN => n1221);
   U1477 : AOI22_X1 port map( A1 => n9518, A2 => n10460, B1 => n9515, B2 => 
                           n10276, ZN => n1222);
   U1478 : OAI221_X1 port map( B1 => n8612, B2 => n9524, C1 => n8580, C2 => 
                           n9521, A => n1204, ZN => n1203);
   U1479 : AOI22_X1 port map( A1 => n9518, A2 => n10459, B1 => n9515, B2 => 
                           n10275, ZN => n1204);
   U1480 : OAI221_X1 port map( B1 => n8613, B2 => n9524, C1 => n8581, C2 => 
                           n9521, A => n1186, ZN => n1185);
   U1481 : AOI22_X1 port map( A1 => n9518, A2 => n10458, B1 => n9515, B2 => 
                           n10274, ZN => n1186);
   U1482 : OAI221_X1 port map( B1 => n2351, B2 => n9487, C1 => n8375, C2 => 
                           n9484, A => n1469, ZN => n1452);
   U1483 : AOI22_X1 port map( A1 => n9481, A2 => n10225, B1 => n9480, B2 => 
                           n10657, ZN => n1469);
   U1484 : OAI221_X1 port map( B1 => n8252, B2 => n9512, C1 => n8218, C2 => 
                           n9509, A => n1223, ZN => n1220);
   U1485 : AOI22_X1 port map( A1 => n9506, A2 => n10596, B1 => n9503, B2 => 
                           n10428, ZN => n1223);
   U1486 : AOI22_X1 port map( A1 => n9434, A2 => n10332, B1 => n9431, B2 => 
                           n9940, ZN => n1233);
   U1487 : AOI22_X1 port map( A1 => n9433, A2 => n10345, B1 => n9432, B2 => 
                           n9953, ZN => n1479);
   U1488 : AOI22_X1 port map( A1 => n9506, A2 => n10595, B1 => n9503, B2 => 
                           n10427, ZN => n1205);
   U1489 : AOI22_X1 port map( A1 => n9506, A2 => n10594, B1 => n9503, B2 => 
                           n10426, ZN => n1187);
   U1490 : AOI22_X1 port map( A1 => n9506, A2 => n10589, B1 => n9502, B2 => 
                           n10421, ZN => n1097);
   U1491 : AOI22_X1 port map( A1 => n9505, A2 => n10599, B1 => n9503, B2 => 
                           n10431, ZN => n1277);
   U1492 : AOI22_X1 port map( A1 => n9505, A2 => n10598, B1 => n9503, B2 => 
                           n10430, ZN => n1259);
   U1493 : AOI22_X1 port map( A1 => n9506, A2 => n10587, B1 => n9502, B2 => 
                           n10419, ZN => n1061);
   U1494 : AOI22_X1 port map( A1 => n9506, A2 => n10588, B1 => n9502, B2 => 
                           n10420, ZN => n1079);
   U1495 : AOI22_X1 port map( A1 => n9506, A2 => n10593, B1 => n9503, B2 => 
                           n10425, ZN => n1169);
   U1496 : AOI22_X1 port map( A1 => n9506, A2 => n10597, B1 => n9503, B2 => 
                           n10429, ZN => n1241);
   U1497 : AOI22_X1 port map( A1 => n9506, A2 => n10586, B1 => n9502, B2 => 
                           n10418, ZN => n1043);
   U1498 : OAI221_X1 port map( B1 => n8615, B2 => n9524, C1 => n8583, C2 => 
                           n9521, A => n1150, ZN => n1149);
   U1499 : AOI22_X1 port map( A1 => n9518, A2 => n10456, B1 => n9515, B2 => 
                           n10272, ZN => n1150);
   U1500 : OAI221_X1 port map( B1 => n8616, B2 => n9524, C1 => n8584, C2 => 
                           n9521, A => n1132, ZN => n1131);
   U1501 : AOI22_X1 port map( A1 => n9518, A2 => n10455, B1 => n9515, B2 => 
                           n10271, ZN => n1132);
   U1502 : OAI221_X1 port map( B1 => n8617, B2 => n9524, C1 => n8585, C2 => 
                           n9521, A => n1114, ZN => n1113);
   U1503 : AOI22_X1 port map( A1 => n9518, A2 => n10454, B1 => n9515, B2 => 
                           n10270, ZN => n1114);
   U1504 : OAI221_X1 port map( B1 => n8256, B2 => n9512, C1 => n8210, C2 => 
                           n9509, A => n1151, ZN => n1148);
   U1505 : AOI22_X1 port map( A1 => n9506, A2 => n10592, B1 => n9503, B2 => 
                           n10424, ZN => n1151);
   U1506 : AOI22_X1 port map( A1 => n9434, A2 => n10328, B1 => n9431, B2 => 
                           n9936, ZN => n1161);
   U1507 : AOI22_X1 port map( A1 => n9506, A2 => n10591, B1 => n9503, B2 => 
                           n10423, ZN => n1133);
   U1508 : AOI22_X1 port map( A1 => n9506, A2 => n10590, B1 => n9503, B2 => 
                           n10422, ZN => n1115);
   U1509 : OAI221_X1 port map( B1 => n2343, B2 => n9487, C1 => n8376, C2 => 
                           n9484, A => n1441, ZN => n1434);
   U1510 : AOI22_X1 port map( A1 => n9481, A2 => n10224, B1 => n9480, B2 => 
                           n10656, ZN => n1441);
   U1511 : AOI22_X1 port map( A1 => n9505, A2 => n10608, B1 => n9504, B2 => 
                           n10440, ZN => n1439);
   U1512 : OAI221_X1 port map( B1 => n8623, B2 => n9525, C1 => n8591, C2 => 
                           n9522, A => n1006, ZN => n1005);
   U1513 : AOI22_X1 port map( A1 => n9519, A2 => n10448, B1 => n9514, B2 => 
                           n10264, ZN => n1006);
   U1514 : OAI221_X1 port map( B1 => n8626, B2 => n9525, C1 => n8594, C2 => 
                           n9522, A => n952, ZN => n951);
   U1515 : AOI22_X1 port map( A1 => n9519, A2 => n10445, B1 => n9514, B2 => 
                           n10261, ZN => n952);
   U1516 : OAI221_X1 port map( B1 => n2335, B2 => n9487, C1 => n8377, C2 => 
                           n9484, A => n1423, ZN => n1416);
   U1517 : AOI22_X1 port map( A1 => n9481, A2 => n10223, B1 => n9480, B2 => 
                           n10655, ZN => n1423);
   U1518 : OAI221_X1 port map( B1 => n2303, B2 => n9487, C1 => n8381, C2 => 
                           n9484, A => n1351, ZN => n1344);
   U1519 : AOI22_X1 port map( A1 => n9481, A2 => n10219, B1 => n9480, B2 => 
                           n10651, ZN => n1351);
   U1520 : OAI221_X1 port map( B1 => n2295, B2 => n9487, C1 => n8382, C2 => 
                           n9484, A => n1333, ZN => n1326);
   U1521 : AOI22_X1 port map( A1 => n9481, A2 => n10218, B1 => n9480, B2 => 
                           n10650, ZN => n1333);
   U1522 : AOI22_X1 port map( A1 => n9505, A2 => n10607, B1 => n9504, B2 => 
                           n10439, ZN => n1421);
   U1523 : AOI22_X1 port map( A1 => n9433, A2 => n10339, B1 => n9432, B2 => 
                           n9947, ZN => n1359);
   U1524 : AOI22_X1 port map( A1 => n9505, A2 => n10602, B1 => n9504, B2 => 
                           n10434, ZN => n1331);
   U1525 : AOI22_X1 port map( A1 => n9505, A2 => n10601, B1 => n9503, B2 => 
                           n10433, ZN => n1313);
   U1526 : AOI22_X1 port map( A1 => n9505, A2 => n10600, B1 => n9503, B2 => 
                           n10432, ZN => n1295);
   U1527 : AOI22_X1 port map( A1 => n9349, A2 => n10041, B1 => n9348, B2 => 
                           n10073, ZN => n2097);
   U1528 : AOI22_X1 port map( A1 => n9361, A2 => n10105, B1 => n9360, B2 => 
                           n10137, ZN => n2096);
   U1529 : AOI22_X1 port map( A1 => n9337, A2 => n9953, B1 => n9336, B2 => 
                           n9985, ZN => n2099);
   U1530 : AOI22_X1 port map( A1 => n9349, A2 => n10040, B1 => n9348, B2 => 
                           n10072, ZN => n2068);
   U1531 : AOI22_X1 port map( A1 => n9361, A2 => n10104, B1 => n9360, B2 => 
                           n10136, ZN => n2067);
   U1532 : AOI22_X1 port map( A1 => n9337, A2 => n9952, B1 => n9336, B2 => 
                           n9984, ZN => n2069);
   U1533 : AOI22_X1 port map( A1 => n9349, A2 => n10039, B1 => n9348, B2 => 
                           n10071, ZN => n2050);
   U1534 : AOI22_X1 port map( A1 => n9361, A2 => n10103, B1 => n9360, B2 => 
                           n10135, ZN => n2049);
   U1535 : AOI22_X1 port map( A1 => n9337, A2 => n9951, B1 => n9336, B2 => 
                           n9983, ZN => n2051);
   U1536 : AOI22_X1 port map( A1 => n9349, A2 => n10038, B1 => n9348, B2 => 
                           n10070, ZN => n2032);
   U1537 : AOI22_X1 port map( A1 => n9361, A2 => n10102, B1 => n9360, B2 => 
                           n10134, ZN => n2031);
   U1538 : AOI22_X1 port map( A1 => n9337, A2 => n9950, B1 => n9336, B2 => 
                           n9982, ZN => n2033);
   U1539 : AOI22_X1 port map( A1 => n9349, A2 => n10037, B1 => n9348, B2 => 
                           n10069, ZN => n2014);
   U1540 : AOI22_X1 port map( A1 => n9361, A2 => n10101, B1 => n9360, B2 => 
                           n10133, ZN => n2013);
   U1541 : AOI22_X1 port map( A1 => n9337, A2 => n9949, B1 => n9336, B2 => 
                           n9981, ZN => n2015);
   U1542 : AOI22_X1 port map( A1 => n9349, A2 => n10036, B1 => n9348, B2 => 
                           n10068, ZN => n1996);
   U1543 : AOI22_X1 port map( A1 => n9361, A2 => n10100, B1 => n9360, B2 => 
                           n10132, ZN => n1995);
   U1544 : AOI22_X1 port map( A1 => n9337, A2 => n9948, B1 => n9336, B2 => 
                           n9980, ZN => n1997);
   U1545 : AOI22_X1 port map( A1 => n9349, A2 => n10035, B1 => n9348, B2 => 
                           n10067, ZN => n1978);
   U1546 : AOI22_X1 port map( A1 => n9361, A2 => n10099, B1 => n9360, B2 => 
                           n10131, ZN => n1977);
   U1547 : AOI22_X1 port map( A1 => n9337, A2 => n9947, B1 => n9336, B2 => 
                           n9979, ZN => n1979);
   U1548 : AOI22_X1 port map( A1 => n9349, A2 => n10034, B1 => n9348, B2 => 
                           n10066, ZN => n1960);
   U1549 : AOI22_X1 port map( A1 => n9361, A2 => n10098, B1 => n9360, B2 => 
                           n10130, ZN => n1959);
   U1550 : AOI22_X1 port map( A1 => n9337, A2 => n9946, B1 => n9336, B2 => 
                           n9978, ZN => n1961);
   U1551 : AOI22_X1 port map( A1 => n9409, A2 => n10625, B1 => n9407, B2 => 
                           n10601, ZN => n1933);
   U1552 : AOI22_X1 port map( A1 => n9397, A2 => n10369, B1 => n9395, B2 => 
                           n10401, ZN => n1934);
   U1553 : AOI22_X1 port map( A1 => n9385, A2 => n10281, B1 => n9383, B2 => 
                           n10313, ZN => n1935);
   U1554 : AOI22_X1 port map( A1 => n9409, A2 => n10624, B1 => n9407, B2 => 
                           n10600, ZN => n1915);
   U1555 : AOI22_X1 port map( A1 => n9397, A2 => n10368, B1 => n9395, B2 => 
                           n10400, ZN => n1916);
   U1556 : AOI22_X1 port map( A1 => n9385, A2 => n10280, B1 => n9383, B2 => 
                           n10312, ZN => n1917);
   U1557 : AOI22_X1 port map( A1 => n9409, A2 => n10623, B1 => n9407, B2 => 
                           n10599, ZN => n1897);
   U1558 : AOI22_X1 port map( A1 => n9397, A2 => n10367, B1 => n9395, B2 => 
                           n10399, ZN => n1898);
   U1559 : AOI22_X1 port map( A1 => n9385, A2 => n10279, B1 => n9383, B2 => 
                           n10311, ZN => n1899);
   U1560 : AOI22_X1 port map( A1 => n9409, A2 => n10622, B1 => n9407, B2 => 
                           n10598, ZN => n1879);
   U1561 : AOI22_X1 port map( A1 => n9397, A2 => n10366, B1 => n9395, B2 => 
                           n10398, ZN => n1880);
   U1562 : AOI22_X1 port map( A1 => n9385, A2 => n10278, B1 => n9383, B2 => 
                           n10310, ZN => n1881);
   U1563 : AOI22_X1 port map( A1 => n9410, A2 => n10621, B1 => n9407, B2 => 
                           n10597, ZN => n1861);
   U1564 : AOI22_X1 port map( A1 => n9398, A2 => n10365, B1 => n9395, B2 => 
                           n10397, ZN => n1862);
   U1565 : AOI22_X1 port map( A1 => n9386, A2 => n10277, B1 => n9383, B2 => 
                           n10309, ZN => n1863);
   U1566 : AOI22_X1 port map( A1 => n9410, A2 => n10620, B1 => n9407, B2 => 
                           n10596, ZN => n1843);
   U1567 : AOI22_X1 port map( A1 => n9398, A2 => n10364, B1 => n9395, B2 => 
                           n10396, ZN => n1844);
   U1568 : AOI22_X1 port map( A1 => n9386, A2 => n10276, B1 => n9383, B2 => 
                           n10308, ZN => n1845);
   U1569 : AOI22_X1 port map( A1 => n9410, A2 => n10619, B1 => n9407, B2 => 
                           n10595, ZN => n1825);
   U1570 : AOI22_X1 port map( A1 => n9398, A2 => n10363, B1 => n9395, B2 => 
                           n10395, ZN => n1826);
   U1571 : AOI22_X1 port map( A1 => n9386, A2 => n10275, B1 => n9383, B2 => 
                           n10307, ZN => n1827);
   U1572 : AOI22_X1 port map( A1 => n9410, A2 => n10618, B1 => n9407, B2 => 
                           n10594, ZN => n1807);
   U1573 : AOI22_X1 port map( A1 => n9398, A2 => n10362, B1 => n9395, B2 => 
                           n10394, ZN => n1808);
   U1574 : AOI22_X1 port map( A1 => n9386, A2 => n10274, B1 => n9383, B2 => 
                           n10306, ZN => n1809);
   U1575 : AOI22_X1 port map( A1 => n9410, A2 => n10617, B1 => n9407, B2 => 
                           n10593, ZN => n1789);
   U1576 : AOI22_X1 port map( A1 => n9398, A2 => n10361, B1 => n9395, B2 => 
                           n10393, ZN => n1790);
   U1577 : AOI22_X1 port map( A1 => n9386, A2 => n10273, B1 => n9383, B2 => 
                           n10305, ZN => n1791);
   U1578 : AOI22_X1 port map( A1 => n9410, A2 => n10616, B1 => n9407, B2 => 
                           n10592, ZN => n1771);
   U1579 : AOI22_X1 port map( A1 => n9398, A2 => n10360, B1 => n9395, B2 => 
                           n10392, ZN => n1772);
   U1580 : AOI22_X1 port map( A1 => n9386, A2 => n10272, B1 => n9383, B2 => 
                           n10304, ZN => n1773);
   U1581 : AOI22_X1 port map( A1 => n9410, A2 => n10615, B1 => n9407, B2 => 
                           n10591, ZN => n1753);
   U1582 : AOI22_X1 port map( A1 => n9398, A2 => n10359, B1 => n9395, B2 => 
                           n10391, ZN => n1754);
   U1583 : AOI22_X1 port map( A1 => n9386, A2 => n10271, B1 => n9383, B2 => 
                           n10303, ZN => n1755);
   U1584 : AOI22_X1 port map( A1 => n9410, A2 => n10614, B1 => n9407, B2 => 
                           n10590, ZN => n1735);
   U1585 : AOI22_X1 port map( A1 => n9398, A2 => n10358, B1 => n9395, B2 => 
                           n10390, ZN => n1736);
   U1586 : AOI22_X1 port map( A1 => n9386, A2 => n10270, B1 => n9383, B2 => 
                           n10302, ZN => n1737);
   U1587 : AOI22_X1 port map( A1 => n9410, A2 => n10613, B1 => n9406, B2 => 
                           n10589, ZN => n1717);
   U1588 : AOI22_X1 port map( A1 => n9398, A2 => n10357, B1 => n9394, B2 => 
                           n10389, ZN => n1718);
   U1589 : AOI22_X1 port map( A1 => n9386, A2 => n10269, B1 => n9382, B2 => 
                           n10301, ZN => n1719);
   U1590 : AOI22_X1 port map( A1 => n9410, A2 => n10612, B1 => n9406, B2 => 
                           n10588, ZN => n1699);
   U1591 : AOI22_X1 port map( A1 => n9398, A2 => n10356, B1 => n9394, B2 => 
                           n10388, ZN => n1700);
   U1592 : AOI22_X1 port map( A1 => n9386, A2 => n10268, B1 => n9382, B2 => 
                           n10300, ZN => n1701);
   U1593 : AOI22_X1 port map( A1 => n9410, A2 => n10611, B1 => n9406, B2 => 
                           n10587, ZN => n1681);
   U1594 : AOI22_X1 port map( A1 => n9398, A2 => n10355, B1 => n9394, B2 => 
                           n10387, ZN => n1682);
   U1595 : AOI22_X1 port map( A1 => n9386, A2 => n10267, B1 => n9382, B2 => 
                           n10299, ZN => n1683);
   U1596 : AOI22_X1 port map( A1 => n9410, A2 => n10610, B1 => n9406, B2 => 
                           n10586, ZN => n1663);
   U1597 : AOI22_X1 port map( A1 => n9398, A2 => n10354, B1 => n9394, B2 => 
                           n10386, ZN => n1664);
   U1598 : AOI22_X1 port map( A1 => n9386, A2 => n10266, B1 => n9382, B2 => 
                           n10298, ZN => n1665);
   U1599 : AOI22_X1 port map( A1 => n9411, A2 => n10553, B1 => n9406, B2 => 
                           n10545, ZN => n1645);
   U1600 : AOI22_X1 port map( A1 => n9399, A2 => n10353, B1 => n9394, B2 => 
                           n10385, ZN => n1646);
   U1601 : AOI22_X1 port map( A1 => n9387, A2 => n10265, B1 => n9382, B2 => 
                           n10297, ZN => n1647);
   U1602 : AOI22_X1 port map( A1 => n9411, A2 => n10552, B1 => n9406, B2 => 
                           n10544, ZN => n1627);
   U1603 : AOI22_X1 port map( A1 => n9399, A2 => n10352, B1 => n9394, B2 => 
                           n10384, ZN => n1628);
   U1604 : AOI22_X1 port map( A1 => n9387, A2 => n10264, B1 => n9382, B2 => 
                           n10296, ZN => n1629);
   U1605 : AOI22_X1 port map( A1 => n9411, A2 => n10551, B1 => n9406, B2 => 
                           n10543, ZN => n1609);
   U1606 : AOI22_X1 port map( A1 => n9399, A2 => n10351, B1 => n9394, B2 => 
                           n10383, ZN => n1610);
   U1607 : AOI22_X1 port map( A1 => n9387, A2 => n10263, B1 => n9382, B2 => 
                           n10295, ZN => n1611);
   U1608 : AOI22_X1 port map( A1 => n9411, A2 => n10550, B1 => n9406, B2 => 
                           n10542, ZN => n1591);
   U1609 : AOI22_X1 port map( A1 => n9399, A2 => n10350, B1 => n9394, B2 => 
                           n10382, ZN => n1592);
   U1610 : AOI22_X1 port map( A1 => n9387, A2 => n10262, B1 => n9382, B2 => 
                           n10294, ZN => n1593);
   U1611 : AOI22_X1 port map( A1 => n9411, A2 => n10549, B1 => n9406, B2 => 
                           n10541, ZN => n1573);
   U1612 : AOI22_X1 port map( A1 => n9399, A2 => n10349, B1 => n9394, B2 => 
                           n10381, ZN => n1574);
   U1613 : AOI22_X1 port map( A1 => n9387, A2 => n10261, B1 => n9382, B2 => 
                           n10293, ZN => n1575);
   U1614 : AOI22_X1 port map( A1 => n9411, A2 => n10548, B1 => n9406, B2 => 
                           n10540, ZN => n1555);
   U1615 : AOI22_X1 port map( A1 => n9399, A2 => n10348, B1 => n9394, B2 => 
                           n10380, ZN => n1556);
   U1616 : AOI22_X1 port map( A1 => n9387, A2 => n10260, B1 => n9382, B2 => 
                           n10292, ZN => n1557);
   U1617 : AOI22_X1 port map( A1 => n9411, A2 => n10547, B1 => n9406, B2 => 
                           n10539, ZN => n1537);
   U1618 : AOI22_X1 port map( A1 => n9399, A2 => n10347, B1 => n9394, B2 => 
                           n10379, ZN => n1538);
   U1619 : AOI22_X1 port map( A1 => n9387, A2 => n10259, B1 => n9382, B2 => 
                           n10291, ZN => n1539);
   U1620 : AOI22_X1 port map( A1 => n9411, A2 => n10546, B1 => n9406, B2 => 
                           n10538, ZN => n1493);
   U1621 : AOI22_X1 port map( A1 => n9399, A2 => n10346, B1 => n9394, B2 => 
                           n10378, ZN => n1498);
   U1622 : AOI22_X1 port map( A1 => n9387, A2 => n10258, B1 => n9382, B2 => 
                           n10290, ZN => n1503);
   U1623 : OAI221_X1 port map( B1 => n8654, B2 => n9379, C1 => n8630, C2 => 
                           n9376, A => n2094, ZN => n2093);
   U1624 : AOI22_X1 port map( A1 => n9373, A2 => n10225, B1 => n9372, B2 => 
                           n10257, ZN => n2094);
   U1625 : OAI221_X1 port map( B1 => n8375, B2 => n9427, C1 => n8343, C2 => 
                           n9424, A => n2076, ZN => n2075);
   U1626 : AOI22_X1 port map( A1 => n9421, A2 => n10657, B1 => n9420, B2 => 
                           n10537, ZN => n2076);
   U1627 : OAI221_X1 port map( B1 => n8439, B2 => n9415, C1 => n8407, C2 => 
                           n9412, A => n2082, ZN => n2074);
   U1628 : AOI22_X1 port map( A1 => n9409, A2 => n10633, B1 => n9408, B2 => 
                           n10609, ZN => n2082);
   U1629 : OAI221_X1 port map( B1 => n8478, B2 => n9403, C1 => n8471, C2 => 
                           n9400, A => n2087, ZN => n2073);
   U1630 : AOI22_X1 port map( A1 => n9397, A2 => n10377, B1 => n9396, B2 => 
                           n10409, ZN => n2087);
   U1631 : OAI221_X1 port map( B1 => n8566, B2 => n9391, C1 => n8542, C2 => 
                           n9388, A => n2089, ZN => n2072);
   U1632 : AOI22_X1 port map( A1 => n9385, A2 => n10289, B1 => n9384, B2 => 
                           n10321, ZN => n2089);
   U1633 : OAI221_X1 port map( B1 => n8655, B2 => n9379, C1 => n8631, C2 => 
                           n9376, A => n2066, ZN => n2065);
   U1634 : AOI22_X1 port map( A1 => n9373, A2 => n10224, B1 => n9372, B2 => 
                           n10256, ZN => n2066);
   U1635 : OAI221_X1 port map( B1 => n8376, B2 => n9427, C1 => n8344, C2 => 
                           n9424, A => n2058, ZN => n2057);
   U1636 : AOI22_X1 port map( A1 => n9421, A2 => n10656, B1 => n9420, B2 => 
                           n10536, ZN => n2058);
   U1637 : OAI221_X1 port map( B1 => n8440, B2 => n9415, C1 => n8408, C2 => 
                           n9412, A => n2059, ZN => n2056);
   U1638 : AOI22_X1 port map( A1 => n9409, A2 => n10632, B1 => n9408, B2 => 
                           n10608, ZN => n2059);
   U1639 : OAI221_X1 port map( B1 => n8479, B2 => n9403, C1 => n8472, C2 => 
                           n9400, A => n2060, ZN => n2055);
   U1640 : AOI22_X1 port map( A1 => n9397, A2 => n10376, B1 => n9396, B2 => 
                           n10408, ZN => n2060);
   U1641 : OAI221_X1 port map( B1 => n8567, B2 => n9391, C1 => n8543, C2 => 
                           n9388, A => n2061, ZN => n2054);
   U1642 : AOI22_X1 port map( A1 => n9385, A2 => n10288, B1 => n9384, B2 => 
                           n10320, ZN => n2061);
   U1643 : OAI221_X1 port map( B1 => n8656, B2 => n9379, C1 => n8632, C2 => 
                           n9376, A => n2048, ZN => n2047);
   U1644 : AOI22_X1 port map( A1 => n9373, A2 => n10223, B1 => n9372, B2 => 
                           n10255, ZN => n2048);
   U1645 : OAI221_X1 port map( B1 => n8377, B2 => n9427, C1 => n8345, C2 => 
                           n9424, A => n2040, ZN => n2039);
   U1646 : AOI22_X1 port map( A1 => n9421, A2 => n10655, B1 => n9420, B2 => 
                           n10535, ZN => n2040);
   U1647 : OAI221_X1 port map( B1 => n8441, B2 => n9415, C1 => n8409, C2 => 
                           n9412, A => n2041, ZN => n2038);
   U1648 : AOI22_X1 port map( A1 => n9409, A2 => n10631, B1 => n9408, B2 => 
                           n10607, ZN => n2041);
   U1649 : OAI221_X1 port map( B1 => n8480, B2 => n9403, C1 => n8473, C2 => 
                           n9400, A => n2042, ZN => n2037);
   U1650 : AOI22_X1 port map( A1 => n9397, A2 => n10375, B1 => n9396, B2 => 
                           n10407, ZN => n2042);
   U1651 : OAI221_X1 port map( B1 => n8568, B2 => n9391, C1 => n8544, C2 => 
                           n9388, A => n2043, ZN => n2036);
   U1652 : AOI22_X1 port map( A1 => n9385, A2 => n10287, B1 => n9384, B2 => 
                           n10319, ZN => n2043);
   U1653 : OAI221_X1 port map( B1 => n8657, B2 => n9379, C1 => n8633, C2 => 
                           n9376, A => n2030, ZN => n2029);
   U1654 : AOI22_X1 port map( A1 => n9373, A2 => n10222, B1 => n9372, B2 => 
                           n10254, ZN => n2030);
   U1655 : OAI221_X1 port map( B1 => n8378, B2 => n9427, C1 => n8346, C2 => 
                           n9424, A => n2022, ZN => n2021);
   U1656 : AOI22_X1 port map( A1 => n9421, A2 => n10654, B1 => n9420, B2 => 
                           n10534, ZN => n2022);
   U1657 : OAI221_X1 port map( B1 => n8442, B2 => n9415, C1 => n8410, C2 => 
                           n9412, A => n2023, ZN => n2020);
   U1658 : AOI22_X1 port map( A1 => n9409, A2 => n10630, B1 => n9408, B2 => 
                           n10606, ZN => n2023);
   U1659 : OAI221_X1 port map( B1 => n8481, B2 => n9403, C1 => n8474, C2 => 
                           n9400, A => n2024, ZN => n2019);
   U1660 : AOI22_X1 port map( A1 => n9397, A2 => n10374, B1 => n9396, B2 => 
                           n10406, ZN => n2024);
   U1661 : OAI221_X1 port map( B1 => n8569, B2 => n9391, C1 => n8545, C2 => 
                           n9388, A => n2025, ZN => n2018);
   U1662 : AOI22_X1 port map( A1 => n9385, A2 => n10286, B1 => n9384, B2 => 
                           n10318, ZN => n2025);
   U1663 : OAI221_X1 port map( B1 => n8658, B2 => n9379, C1 => n8634, C2 => 
                           n9376, A => n2012, ZN => n2011);
   U1664 : AOI22_X1 port map( A1 => n9373, A2 => n10221, B1 => n9372, B2 => 
                           n10253, ZN => n2012);
   U1665 : OAI221_X1 port map( B1 => n8379, B2 => n9427, C1 => n8347, C2 => 
                           n9424, A => n2004, ZN => n2003);
   U1666 : AOI22_X1 port map( A1 => n9421, A2 => n10653, B1 => n9420, B2 => 
                           n10533, ZN => n2004);
   U1667 : OAI221_X1 port map( B1 => n8443, B2 => n9415, C1 => n8411, C2 => 
                           n9412, A => n2005, ZN => n2002);
   U1668 : AOI22_X1 port map( A1 => n9409, A2 => n10629, B1 => n9408, B2 => 
                           n10605, ZN => n2005);
   U1669 : OAI221_X1 port map( B1 => n8482, B2 => n9403, C1 => n8475, C2 => 
                           n9400, A => n2006, ZN => n2001);
   U1670 : AOI22_X1 port map( A1 => n9397, A2 => n10373, B1 => n9396, B2 => 
                           n10405, ZN => n2006);
   U1671 : OAI221_X1 port map( B1 => n8570, B2 => n9391, C1 => n8546, C2 => 
                           n9388, A => n2007, ZN => n2000);
   U1672 : AOI22_X1 port map( A1 => n9385, A2 => n10285, B1 => n9384, B2 => 
                           n10317, ZN => n2007);
   U1673 : OAI221_X1 port map( B1 => n8659, B2 => n9379, C1 => n8635, C2 => 
                           n9376, A => n1994, ZN => n1993);
   U1674 : AOI22_X1 port map( A1 => n9373, A2 => n10220, B1 => n9372, B2 => 
                           n10252, ZN => n1994);
   U1675 : OAI221_X1 port map( B1 => n8380, B2 => n9427, C1 => n8348, C2 => 
                           n9424, A => n1986, ZN => n1985);
   U1676 : AOI22_X1 port map( A1 => n9421, A2 => n10652, B1 => n9420, B2 => 
                           n10532, ZN => n1986);
   U1677 : OAI221_X1 port map( B1 => n8444, B2 => n9415, C1 => n8412, C2 => 
                           n9412, A => n1987, ZN => n1984);
   U1678 : AOI22_X1 port map( A1 => n9409, A2 => n10628, B1 => n9408, B2 => 
                           n10604, ZN => n1987);
   U1679 : OAI221_X1 port map( B1 => n8483, B2 => n9403, C1 => n8476, C2 => 
                           n9400, A => n1988, ZN => n1983);
   U1680 : AOI22_X1 port map( A1 => n9397, A2 => n10372, B1 => n9396, B2 => 
                           n10404, ZN => n1988);
   U1681 : OAI221_X1 port map( B1 => n8571, B2 => n9391, C1 => n8547, C2 => 
                           n9388, A => n1989, ZN => n1982);
   U1682 : AOI22_X1 port map( A1 => n9385, A2 => n10284, B1 => n9384, B2 => 
                           n10316, ZN => n1989);
   U1683 : OAI221_X1 port map( B1 => n8660, B2 => n9379, C1 => n8636, C2 => 
                           n9376, A => n1976, ZN => n1975);
   U1684 : AOI22_X1 port map( A1 => n9373, A2 => n10219, B1 => n9372, B2 => 
                           n10251, ZN => n1976);
   U1685 : OAI221_X1 port map( B1 => n8381, B2 => n9427, C1 => n8349, C2 => 
                           n9424, A => n1968, ZN => n1967);
   U1687 : AOI22_X1 port map( A1 => n9421, A2 => n10651, B1 => n9420, B2 => 
                           n10531, ZN => n1968);
   U1688 : OAI221_X1 port map( B1 => n8445, B2 => n9415, C1 => n8413, C2 => 
                           n9412, A => n1969, ZN => n1966);
   U1689 : AOI22_X1 port map( A1 => n9409, A2 => n10627, B1 => n9408, B2 => 
                           n10603, ZN => n1969);
   U1690 : OAI221_X1 port map( B1 => n8484, B2 => n9403, C1 => n8477, C2 => 
                           n9400, A => n1970, ZN => n1965);
   U1691 : AOI22_X1 port map( A1 => n9397, A2 => n10371, B1 => n9396, B2 => 
                           n10403, ZN => n1970);
   U1692 : OAI221_X1 port map( B1 => n8572, B2 => n9391, C1 => n8548, C2 => 
                           n9388, A => n1971, ZN => n1964);
   U1693 : AOI22_X1 port map( A1 => n9385, A2 => n10283, B1 => n9384, B2 => 
                           n10315, ZN => n1971);
   U1694 : OAI221_X1 port map( B1 => n8661, B2 => n9379, C1 => n8637, C2 => 
                           n9376, A => n1958, ZN => n1957);
   U1695 : AOI22_X1 port map( A1 => n9373, A2 => n10218, B1 => n9372, B2 => 
                           n10250, ZN => n1958);
   U1696 : OAI221_X1 port map( B1 => n8382, B2 => n9427, C1 => n8350, C2 => 
                           n9424, A => n1950, ZN => n1949);
   U1697 : AOI22_X1 port map( A1 => n9421, A2 => n10650, B1 => n9420, B2 => 
                           n10530, ZN => n1950);
   U1698 : OAI221_X1 port map( B1 => n8446, B2 => n9415, C1 => n8414, C2 => 
                           n9412, A => n1951, ZN => n1948);
   U1700 : AOI22_X1 port map( A1 => n9409, A2 => n10626, B1 => n9408, B2 => 
                           n10602, ZN => n1951);
   U1701 : OAI221_X1 port map( B1 => n8485, B2 => n9403, C1 => n8246, C2 => 
                           n9400, A => n1952, ZN => n1947);
   U1702 : AOI22_X1 port map( A1 => n9397, A2 => n10370, B1 => n9396, B2 => 
                           n10402, ZN => n1952);
   U1703 : OAI221_X1 port map( B1 => n8573, B2 => n9391, C1 => n8549, C2 => 
                           n9388, A => n1953, ZN => n1946);
   U1704 : AOI22_X1 port map( A1 => n9385, A2 => n10282, B1 => n9384, B2 => 
                           n10314, ZN => n1953);
   U1705 : OAI221_X1 port map( B1 => n8383, B2 => n9427, C1 => n8351, C2 => 
                           n9424, A => n1932, ZN => n1931);
   U1706 : AOI22_X1 port map( A1 => n9421, A2 => n10649, B1 => n9419, B2 => 
                           n10529, ZN => n1932);
   U1707 : OAI221_X1 port map( B1 => n8750, B2 => n9367, C1 => n8726, C2 => 
                           n9364, A => n1941, ZN => n1938);
   U1708 : AOI22_X1 port map( A1 => n9361, A2 => n10097, B1 => n9359, B2 => 
                           n10129, ZN => n1941);
   U1709 : OAI221_X1 port map( B1 => n8384, B2 => n9427, C1 => n8352, C2 => 
                           n9424, A => n1914, ZN => n1913);
   U1710 : AOI22_X1 port map( A1 => n9421, A2 => n10648, B1 => n9419, B2 => 
                           n10528, ZN => n1914);
   U1711 : OAI221_X1 port map( B1 => n8751, B2 => n9367, C1 => n8727, C2 => 
                           n9364, A => n1923, ZN => n1920);
   U1712 : AOI22_X1 port map( A1 => n9361, A2 => n10096, B1 => n9359, B2 => 
                           n10128, ZN => n1923);
   U1713 : OAI221_X1 port map( B1 => n8385, B2 => n9427, C1 => n8353, C2 => 
                           n9424, A => n1896, ZN => n1895);
   U1714 : AOI22_X1 port map( A1 => n9421, A2 => n10647, B1 => n9419, B2 => 
                           n10527, ZN => n1896);
   U1715 : OAI221_X1 port map( B1 => n8752, B2 => n9367, C1 => n8728, C2 => 
                           n9364, A => n1905, ZN => n1902);
   U1717 : AOI22_X1 port map( A1 => n9361, A2 => n10095, B1 => n9359, B2 => 
                           n10127, ZN => n1905);
   U1718 : OAI221_X1 port map( B1 => n8386, B2 => n9427, C1 => n8354, C2 => 
                           n9424, A => n1878, ZN => n1877);
   U1719 : AOI22_X1 port map( A1 => n9421, A2 => n10646, B1 => n9419, B2 => 
                           n10526, ZN => n1878);
   U1720 : OAI221_X1 port map( B1 => n8753, B2 => n9367, C1 => n8729, C2 => 
                           n9364, A => n1887, ZN => n1884);
   U1721 : AOI22_X1 port map( A1 => n9361, A2 => n10094, B1 => n9359, B2 => 
                           n10126, ZN => n1887);
   U1723 : OAI221_X1 port map( B1 => n8387, B2 => n9428, C1 => n8355, C2 => 
                           n9425, A => n1860, ZN => n1859);
   U1724 : AOI22_X1 port map( A1 => n9422, A2 => n10645, B1 => n9419, B2 => 
                           n10525, ZN => n1860);
   U1725 : OAI221_X1 port map( B1 => n8754, B2 => n9368, C1 => n8730, C2 => 
                           n9365, A => n1869, ZN => n1866);
   U1726 : AOI22_X1 port map( A1 => n9362, A2 => n10093, B1 => n9359, B2 => 
                           n10125, ZN => n1869);
   U1727 : OAI221_X1 port map( B1 => n8388, B2 => n9428, C1 => n8356, C2 => 
                           n9425, A => n1842, ZN => n1841);
   U1728 : AOI22_X1 port map( A1 => n9422, A2 => n10644, B1 => n9419, B2 => 
                           n10524, ZN => n1842);
   U1729 : OAI221_X1 port map( B1 => n8755, B2 => n9368, C1 => n8731, C2 => 
                           n9365, A => n1851, ZN => n1848);
   U1730 : AOI22_X1 port map( A1 => n9362, A2 => n10092, B1 => n9359, B2 => 
                           n10124, ZN => n1851);
   U1731 : OAI221_X1 port map( B1 => n8389, B2 => n9428, C1 => n8357, C2 => 
                           n9425, A => n1824, ZN => n1823);
   U1732 : AOI22_X1 port map( A1 => n9422, A2 => n10643, B1 => n9419, B2 => 
                           n10523, ZN => n1824);
   U1733 : OAI221_X1 port map( B1 => n8756, B2 => n9368, C1 => n8732, C2 => 
                           n9365, A => n1833, ZN => n1830);
   U1734 : AOI22_X1 port map( A1 => n9362, A2 => n10091, B1 => n9359, B2 => 
                           n10123, ZN => n1833);
   U1735 : OAI221_X1 port map( B1 => n8390, B2 => n9428, C1 => n8358, C2 => 
                           n9425, A => n1806, ZN => n1805);
   U1736 : AOI22_X1 port map( A1 => n9422, A2 => n10642, B1 => n9419, B2 => 
                           n10522, ZN => n1806);
   U1737 : OAI221_X1 port map( B1 => n8757, B2 => n9368, C1 => n8733, C2 => 
                           n9365, A => n1815, ZN => n1812);
   U1738 : AOI22_X1 port map( A1 => n9362, A2 => n10090, B1 => n9359, B2 => 
                           n10122, ZN => n1815);
   U1739 : OAI221_X1 port map( B1 => n8391, B2 => n9428, C1 => n8359, C2 => 
                           n9425, A => n1788, ZN => n1787);
   U1740 : AOI22_X1 port map( A1 => n9422, A2 => n10641, B1 => n9419, B2 => 
                           n10521, ZN => n1788);
   U1741 : OAI221_X1 port map( B1 => n8758, B2 => n9368, C1 => n8734, C2 => 
                           n9365, A => n1797, ZN => n1794);
   U1742 : AOI22_X1 port map( A1 => n9362, A2 => n10089, B1 => n9359, B2 => 
                           n10121, ZN => n1797);
   U1743 : OAI221_X1 port map( B1 => n8392, B2 => n9428, C1 => n8360, C2 => 
                           n9425, A => n1770, ZN => n1769);
   U1744 : AOI22_X1 port map( A1 => n9422, A2 => n10640, B1 => n9419, B2 => 
                           n10520, ZN => n1770);
   U1745 : OAI221_X1 port map( B1 => n8759, B2 => n9368, C1 => n8735, C2 => 
                           n9365, A => n1779, ZN => n1776);
   U1746 : AOI22_X1 port map( A1 => n9362, A2 => n10088, B1 => n9359, B2 => 
                           n10120, ZN => n1779);
   U1747 : OAI221_X1 port map( B1 => n8393, B2 => n9428, C1 => n8361, C2 => 
                           n9425, A => n1752, ZN => n1751);
   U1748 : AOI22_X1 port map( A1 => n9422, A2 => n10639, B1 => n9419, B2 => 
                           n10519, ZN => n1752);
   U1749 : OAI221_X1 port map( B1 => n8760, B2 => n9368, C1 => n8736, C2 => 
                           n9365, A => n1761, ZN => n1758);
   U1750 : AOI22_X1 port map( A1 => n9362, A2 => n10087, B1 => n9359, B2 => 
                           n10119, ZN => n1761);
   U1751 : OAI221_X1 port map( B1 => n8394, B2 => n9428, C1 => n8362, C2 => 
                           n9425, A => n1734, ZN => n1733);
   U1752 : AOI22_X1 port map( A1 => n9422, A2 => n10638, B1 => n9419, B2 => 
                           n10518, ZN => n1734);
   U1753 : OAI221_X1 port map( B1 => n8761, B2 => n9368, C1 => n8737, C2 => 
                           n9365, A => n1743, ZN => n1740);
   U1754 : AOI22_X1 port map( A1 => n9362, A2 => n10086, B1 => n9359, B2 => 
                           n10118, ZN => n1743);
   U1755 : OAI221_X1 port map( B1 => n8395, B2 => n9428, C1 => n8363, C2 => 
                           n9425, A => n1716, ZN => n1715);
   U1756 : AOI22_X1 port map( A1 => n9422, A2 => n10637, B1 => n9418, B2 => 
                           n10517, ZN => n1716);
   U1757 : OAI221_X1 port map( B1 => n8762, B2 => n9368, C1 => n8738, C2 => 
                           n9365, A => n1725, ZN => n1722);
   U1758 : AOI22_X1 port map( A1 => n9362, A2 => n10085, B1 => n9358, B2 => 
                           n10117, ZN => n1725);
   U1759 : OAI221_X1 port map( B1 => n8396, B2 => n9428, C1 => n8364, C2 => 
                           n9425, A => n1698, ZN => n1697);
   U1760 : AOI22_X1 port map( A1 => n9422, A2 => n10636, B1 => n9418, B2 => 
                           n10516, ZN => n1698);
   U1761 : OAI221_X1 port map( B1 => n8763, B2 => n9368, C1 => n8739, C2 => 
                           n9365, A => n1707, ZN => n1704);
   U1762 : AOI22_X1 port map( A1 => n9362, A2 => n10084, B1 => n9358, B2 => 
                           n10116, ZN => n1707);
   U1763 : OAI221_X1 port map( B1 => n8397, B2 => n9428, C1 => n8365, C2 => 
                           n9425, A => n1680, ZN => n1679);
   U1764 : AOI22_X1 port map( A1 => n9422, A2 => n10635, B1 => n9418, B2 => 
                           n10515, ZN => n1680);
   U1765 : OAI221_X1 port map( B1 => n8764, B2 => n9368, C1 => n8740, C2 => 
                           n9365, A => n1689, ZN => n1686);
   U1766 : AOI22_X1 port map( A1 => n9362, A2 => n10083, B1 => n9358, B2 => 
                           n10115, ZN => n1689);
   U1767 : OAI221_X1 port map( B1 => n8398, B2 => n9428, C1 => n8366, C2 => 
                           n9425, A => n1662, ZN => n1661);
   U1768 : AOI22_X1 port map( A1 => n9422, A2 => n10634, B1 => n9418, B2 => 
                           n10514, ZN => n1662);
   U1769 : OAI221_X1 port map( B1 => n8765, B2 => n9368, C1 => n8741, C2 => 
                           n9365, A => n1671, ZN => n1668);
   U1770 : AOI22_X1 port map( A1 => n9362, A2 => n10082, B1 => n9358, B2 => 
                           n10114, ZN => n1671);
   U1771 : OAI221_X1 port map( B1 => n8399, B2 => n9429, C1 => n8367, C2 => 
                           n9426, A => n1644, ZN => n1643);
   U1772 : AOI22_X1 port map( A1 => n9423, A2 => n10561, B1 => n9418, B2 => 
                           n10513, ZN => n1644);
   U1773 : OAI221_X1 port map( B1 => n8766, B2 => n9369, C1 => n8287, C2 => 
                           n9366, A => n1653, ZN => n1650);
   U1774 : AOI22_X1 port map( A1 => n9363, A2 => n10081, B1 => n9358, B2 => 
                           n10113, ZN => n1653);
   U1775 : OAI221_X1 port map( B1 => n8400, B2 => n9429, C1 => n8368, C2 => 
                           n9426, A => n1626, ZN => n1625);
   U1776 : AOI22_X1 port map( A1 => n9423, A2 => n10560, B1 => n9418, B2 => 
                           n10512, ZN => n1626);
   U1777 : OAI221_X1 port map( B1 => n8767, B2 => n9369, C1 => n8288, C2 => 
                           n9366, A => n1635, ZN => n1632);
   U1778 : AOI22_X1 port map( A1 => n9363, A2 => n10080, B1 => n9358, B2 => 
                           n10112, ZN => n1635);
   U1779 : OAI221_X1 port map( B1 => n8401, B2 => n9429, C1 => n8369, C2 => 
                           n9426, A => n1608, ZN => n1607);
   U1780 : AOI22_X1 port map( A1 => n9423, A2 => n10559, B1 => n9418, B2 => 
                           n10511, ZN => n1608);
   U1781 : OAI221_X1 port map( B1 => n8768, B2 => n9369, C1 => n8289, C2 => 
                           n9366, A => n1617, ZN => n1614);
   U1782 : AOI22_X1 port map( A1 => n9363, A2 => n10079, B1 => n9358, B2 => 
                           n10111, ZN => n1617);
   U1783 : OAI221_X1 port map( B1 => n8402, B2 => n9429, C1 => n8370, C2 => 
                           n9426, A => n1590, ZN => n1589);
   U1784 : AOI22_X1 port map( A1 => n9423, A2 => n10558, B1 => n9418, B2 => 
                           n10510, ZN => n1590);
   U1785 : OAI221_X1 port map( B1 => n8769, B2 => n9369, C1 => n8290, C2 => 
                           n9366, A => n1599, ZN => n1596);
   U1786 : AOI22_X1 port map( A1 => n9363, A2 => n10078, B1 => n9358, B2 => 
                           n10110, ZN => n1599);
   U1787 : OAI221_X1 port map( B1 => n8403, B2 => n9429, C1 => n8371, C2 => 
                           n9426, A => n1572, ZN => n1571);
   U1788 : AOI22_X1 port map( A1 => n9423, A2 => n10557, B1 => n9418, B2 => 
                           n10509, ZN => n1572);
   U1789 : OAI221_X1 port map( B1 => n8770, B2 => n9369, C1 => n8291, C2 => 
                           n9366, A => n1581, ZN => n1578);
   U1790 : AOI22_X1 port map( A1 => n9363, A2 => n10077, B1 => n9358, B2 => 
                           n10109, ZN => n1581);
   U1791 : OAI221_X1 port map( B1 => n8404, B2 => n9429, C1 => n8372, C2 => 
                           n9426, A => n1554, ZN => n1553);
   U1792 : AOI22_X1 port map( A1 => n9423, A2 => n10556, B1 => n9418, B2 => 
                           n10508, ZN => n1554);
   U1793 : OAI221_X1 port map( B1 => n8771, B2 => n9369, C1 => n8292, C2 => 
                           n9366, A => n1563, ZN => n1560);
   U1794 : AOI22_X1 port map( A1 => n9363, A2 => n10076, B1 => n9358, B2 => 
                           n10108, ZN => n1563);
   U1795 : OAI221_X1 port map( B1 => n8405, B2 => n9429, C1 => n8373, C2 => 
                           n9426, A => n1536, ZN => n1535);
   U1796 : AOI22_X1 port map( A1 => n9423, A2 => n10555, B1 => n9418, B2 => 
                           n10507, ZN => n1536);
   U1797 : OAI221_X1 port map( B1 => n8772, B2 => n9369, C1 => n8293, C2 => 
                           n9366, A => n1545, ZN => n1542);
   U1798 : AOI22_X1 port map( A1 => n9363, A2 => n10075, B1 => n9358, B2 => 
                           n10107, ZN => n1545);
   U1799 : OAI221_X1 port map( B1 => n8406, B2 => n9429, C1 => n8374, C2 => 
                           n9426, A => n1488, ZN => n1485);
   U1800 : AOI22_X1 port map( A1 => n9423, A2 => n10554, B1 => n9418, B2 => 
                           n10506, ZN => n1488);
   U1801 : OAI221_X1 port map( B1 => n8773, B2 => n9369, C1 => n8294, C2 => 
                           n9366, A => n1517, ZN => n1508);
   U1802 : AOI22_X1 port map( A1 => n9363, A2 => n10074, B1 => n9358, B2 => 
                           n10106, ZN => n1517);
   U1803 : OAI22_X1 port map( A1 => n9329, A2 => n9603, B1 => n8655, B2 => 
                           n9612, ZN => n3199);
   U1804 : OAI22_X1 port map( A1 => n9326, A2 => n9603, B1 => n8656, B2 => 
                           n9612, ZN => n3200);
   U1805 : OAI22_X1 port map( A1 => n9323, A2 => n9603, B1 => n8657, B2 => 
                           n9612, ZN => n3201);
   U1806 : OAI22_X1 port map( A1 => n9320, A2 => n9603, B1 => n8658, B2 => 
                           n9611, ZN => n3202);
   U1807 : OAI22_X1 port map( A1 => n9317, A2 => n9603, B1 => n8659, B2 => 
                           n9611, ZN => n3203);
   U1808 : OAI22_X1 port map( A1 => n9311, A2 => n9603, B1 => n8661, B2 => 
                           n9611, ZN => n3205);
   U1809 : OAI22_X1 port map( A1 => n9308, A2 => n9603, B1 => n8662, B2 => 
                           n9610, ZN => n3206);
   U1810 : OAI22_X1 port map( A1 => n9305, A2 => n9603, B1 => n8663, B2 => 
                           n9610, ZN => n3207);
   U1811 : OAI22_X1 port map( A1 => n9302, A2 => n9603, B1 => n8664, B2 => 
                           n9610, ZN => n3208);
   U1812 : OAI22_X1 port map( A1 => n9299, A2 => n9603, B1 => n8665, B2 => 
                           n9610, ZN => n3209);
   U1813 : OAI22_X1 port map( A1 => n9296, A2 => n9604, B1 => n8666, B2 => 
                           n9609, ZN => n3210);
   U1814 : OAI22_X1 port map( A1 => n9290, A2 => n9604, B1 => n8668, B2 => 
                           n9609, ZN => n3212);
   U1815 : OAI22_X1 port map( A1 => n9287, A2 => n9604, B1 => n8669, B2 => 
                           n9609, ZN => n3213);
   U1816 : OAI22_X1 port map( A1 => n9284, A2 => n9604, B1 => n8670, B2 => 
                           n9608, ZN => n3214);
   U1817 : OAI22_X1 port map( A1 => n9278, A2 => n9604, B1 => n8672, B2 => 
                           n9608, ZN => n3216);
   U1818 : OAI22_X1 port map( A1 => n9275, A2 => n9604, B1 => n8673, B2 => 
                           n9608, ZN => n3217);
   U1819 : OAI22_X1 port map( A1 => n9272, A2 => n9604, B1 => n8674, B2 => 
                           n9607, ZN => n3218);
   U1820 : OAI22_X1 port map( A1 => n9269, A2 => n9604, B1 => n8675, B2 => 
                           n9607, ZN => n3219);
   U1821 : OAI22_X1 port map( A1 => n9266, A2 => n9604, B1 => n8676, B2 => 
                           n9607, ZN => n3220);
   U1822 : OAI22_X1 port map( A1 => n9263, A2 => n9604, B1 => n8677, B2 => 
                           n9607, ZN => n3221);
   U1823 : OAI22_X1 port map( A1 => n9260, A2 => n9603, B1 => n8678, B2 => 
                           n9606, ZN => n3222);
   U1824 : OAI22_X1 port map( A1 => n9257, A2 => n9604, B1 => n8679, B2 => 
                           n9606, ZN => n3223);
   U1825 : OAI22_X1 port map( A1 => n9254, A2 => n9603, B1 => n8680, B2 => 
                           n9606, ZN => n3224);
   U1826 : OAI22_X1 port map( A1 => n9251, A2 => n9604, B1 => n8681, B2 => 
                           n9606, ZN => n3225);
   U1827 : OAI22_X1 port map( A1 => n9248, A2 => n9603, B1 => n8682, B2 => 
                           n9605, ZN => n3226);
   U1828 : OAI22_X1 port map( A1 => n9245, A2 => n9604, B1 => n8683, B2 => 
                           n9605, ZN => n3227);
   U1829 : OAI22_X1 port map( A1 => n9242, A2 => n9603, B1 => n8684, B2 => 
                           n9605, ZN => n3228);
   U1830 : OAI22_X1 port map( A1 => n9239, A2 => n9604, B1 => n8685, B2 => 
                           n9605, ZN => n3229);
   U1831 : OAI22_X1 port map( A1 => n9331, A2 => n9835, B1 => n2351, B2 => 
                           n9836, ZN => n9109);
   U1832 : OAI22_X1 port map( A1 => n9328, A2 => n9834, B1 => n2343, B2 => 
                           n9836, ZN => n9108);
   U1833 : OAI22_X1 port map( A1 => n9325, A2 => n9835, B1 => n2335, B2 => 
                           n9836, ZN => n9107);
   U1834 : OAI22_X1 port map( A1 => n9322, A2 => n9834, B1 => n2327, B2 => 
                           n9836, ZN => n9106);
   U1835 : OAI22_X1 port map( A1 => n9319, A2 => n9835, B1 => n2319, B2 => 
                           n9837, ZN => n9105);
   U1836 : OAI22_X1 port map( A1 => n9316, A2 => n9834, B1 => n2311, B2 => 
                           n9837, ZN => n9104);
   U1837 : OAI22_X1 port map( A1 => n9313, A2 => n9835, B1 => n2303, B2 => 
                           n9837, ZN => n9103);
   U1838 : OAI22_X1 port map( A1 => n9310, A2 => n9834, B1 => n2295, B2 => 
                           n9837, ZN => n9102);
   U1839 : OAI22_X1 port map( A1 => n9307, A2 => n9835, B1 => n2287, B2 => 
                           n9838, ZN => n9101);
   U1840 : OAI22_X1 port map( A1 => n9304, A2 => n9835, B1 => n2279, B2 => 
                           n9838, ZN => n9100);
   U1841 : OAI22_X1 port map( A1 => n9301, A2 => n9835, B1 => n2271, B2 => 
                           n9838, ZN => n9099);
   U1842 : OAI22_X1 port map( A1 => n9298, A2 => n9835, B1 => n2263, B2 => 
                           n9838, ZN => n9098);
   U1843 : OAI22_X1 port map( A1 => n9295, A2 => n9835, B1 => n2255, B2 => 
                           n9839, ZN => n9097);
   U1844 : OAI22_X1 port map( A1 => n9292, A2 => n9835, B1 => n2247, B2 => 
                           n9839, ZN => n9096);
   U1845 : OAI22_X1 port map( A1 => n9289, A2 => n9835, B1 => n2239, B2 => 
                           n9839, ZN => n9095);
   U1846 : OAI22_X1 port map( A1 => n9286, A2 => n9835, B1 => n2231, B2 => 
                           n9839, ZN => n9094);
   U1847 : OAI22_X1 port map( A1 => n9283, A2 => n9835, B1 => n2223, B2 => 
                           n9840, ZN => n9093);
   U1848 : OAI22_X1 port map( A1 => n9280, A2 => n9835, B1 => n2215, B2 => 
                           n9840, ZN => n9092);
   U1849 : OAI22_X1 port map( A1 => n9277, A2 => n9835, B1 => n2207, B2 => 
                           n9840, ZN => n9091);
   U1850 : OAI22_X1 port map( A1 => n9274, A2 => n9835, B1 => n2199, B2 => 
                           n9840, ZN => n9090);
   U1851 : OAI22_X1 port map( A1 => n9271, A2 => n9834, B1 => n2191, B2 => 
                           n9841, ZN => n9089);
   U1852 : OAI22_X1 port map( A1 => n9268, A2 => n9834, B1 => n2183, B2 => 
                           n9841, ZN => n9088);
   U1853 : OAI22_X1 port map( A1 => n9265, A2 => n9834, B1 => n2175, B2 => 
                           n9841, ZN => n9087);
   U1854 : OAI22_X1 port map( A1 => n9262, A2 => n9834, B1 => n2167, B2 => 
                           n9841, ZN => n9086);
   U1855 : OAI22_X1 port map( A1 => n9259, A2 => n9834, B1 => n2159, B2 => 
                           n9842, ZN => n9085);
   U1856 : OAI22_X1 port map( A1 => n9256, A2 => n9834, B1 => n2151, B2 => 
                           n9842, ZN => n9084);
   U1857 : OAI22_X1 port map( A1 => n9253, A2 => n9834, B1 => n2143, B2 => 
                           n9842, ZN => n9083);
   U1858 : OAI22_X1 port map( A1 => n9250, A2 => n9834, B1 => n2135, B2 => 
                           n9842, ZN => n9082);
   U1859 : OAI22_X1 port map( A1 => n9247, A2 => n9834, B1 => n2127, B2 => 
                           n9843, ZN => n9081);
   U1860 : OAI22_X1 port map( A1 => n9244, A2 => n9834, B1 => n2119, B2 => 
                           n9843, ZN => n9080);
   U1861 : OAI22_X1 port map( A1 => n9241, A2 => n9834, B1 => n2111, B2 => 
                           n9843, ZN => n9079);
   U1862 : OAI22_X1 port map( A1 => n9238, A2 => n9834, B1 => n2103, B2 => 
                           n9843, ZN => n9078);
   U1863 : OAI22_X1 port map( A1 => n9331, A2 => n9747, B1 => n8439, B2 => 
                           n9748, ZN => n3955);
   U1864 : OAI22_X1 port map( A1 => n9328, A2 => n9746, B1 => n8440, B2 => 
                           n9748, ZN => n3939);
   U1865 : OAI22_X1 port map( A1 => n9325, A2 => n9747, B1 => n8441, B2 => 
                           n9748, ZN => n3923);
   U1866 : OAI22_X1 port map( A1 => n9322, A2 => n9746, B1 => n8442, B2 => 
                           n9748, ZN => n3907);
   U1867 : OAI22_X1 port map( A1 => n9319, A2 => n9747, B1 => n8443, B2 => 
                           n9749, ZN => n3891);
   U1868 : OAI22_X1 port map( A1 => n9316, A2 => n9746, B1 => n8444, B2 => 
                           n9749, ZN => n3875);
   U1869 : OAI22_X1 port map( A1 => n9313, A2 => n9747, B1 => n8445, B2 => 
                           n9749, ZN => n3859);
   U1870 : OAI22_X1 port map( A1 => n9310, A2 => n9746, B1 => n8446, B2 => 
                           n9749, ZN => n3843);
   U1871 : OAI22_X1 port map( A1 => n9307, A2 => n9747, B1 => n8447, B2 => 
                           n9750, ZN => n3827);
   U1872 : OAI22_X1 port map( A1 => n9304, A2 => n9747, B1 => n8448, B2 => 
                           n9750, ZN => n3811);
   U1873 : OAI22_X1 port map( A1 => n9301, A2 => n9747, B1 => n8449, B2 => 
                           n9750, ZN => n3795);
   U1874 : OAI22_X1 port map( A1 => n9298, A2 => n9747, B1 => n8450, B2 => 
                           n9750, ZN => n3779);
   U1875 : OAI22_X1 port map( A1 => n9295, A2 => n9747, B1 => n8451, B2 => 
                           n9751, ZN => n3763);
   U1876 : OAI22_X1 port map( A1 => n9292, A2 => n9747, B1 => n8452, B2 => 
                           n9751, ZN => n3747);
   U1877 : OAI22_X1 port map( A1 => n9289, A2 => n9747, B1 => n8453, B2 => 
                           n9751, ZN => n3731);
   U1878 : OAI22_X1 port map( A1 => n9286, A2 => n9747, B1 => n8454, B2 => 
                           n9751, ZN => n3715);
   U1879 : OAI22_X1 port map( A1 => n9283, A2 => n9747, B1 => n8455, B2 => 
                           n9752, ZN => n3699);
   U1880 : OAI22_X1 port map( A1 => n9280, A2 => n9747, B1 => n8456, B2 => 
                           n9752, ZN => n3683);
   U1881 : OAI22_X1 port map( A1 => n9277, A2 => n9747, B1 => n8457, B2 => 
                           n9752, ZN => n3667);
   U1882 : OAI22_X1 port map( A1 => n9274, A2 => n9747, B1 => n8458, B2 => 
                           n9752, ZN => n3651);
   U1883 : OAI22_X1 port map( A1 => n9271, A2 => n9746, B1 => n8459, B2 => 
                           n9753, ZN => n3635);
   U1884 : OAI22_X1 port map( A1 => n9268, A2 => n9746, B1 => n8460, B2 => 
                           n9753, ZN => n3619);
   U1885 : OAI22_X1 port map( A1 => n9265, A2 => n9746, B1 => n8461, B2 => 
                           n9753, ZN => n3603);
   U1886 : OAI22_X1 port map( A1 => n9262, A2 => n9746, B1 => n8462, B2 => 
                           n9753, ZN => n3587);
   U1887 : OAI22_X1 port map( A1 => n9259, A2 => n9746, B1 => n8463, B2 => 
                           n9754, ZN => n3571);
   U1888 : OAI22_X1 port map( A1 => n9256, A2 => n9746, B1 => n8464, B2 => 
                           n9754, ZN => n3555);
   U1889 : OAI22_X1 port map( A1 => n9253, A2 => n9746, B1 => n8465, B2 => 
                           n9754, ZN => n3539);
   U1890 : OAI22_X1 port map( A1 => n9250, A2 => n9746, B1 => n8466, B2 => 
                           n9754, ZN => n3523);
   U1891 : OAI22_X1 port map( A1 => n9247, A2 => n9746, B1 => n8467, B2 => 
                           n9755, ZN => n3507);
   U1892 : OAI22_X1 port map( A1 => n9244, A2 => n9746, B1 => n8468, B2 => 
                           n9755, ZN => n3491);
   U1893 : OAI22_X1 port map( A1 => n9241, A2 => n9746, B1 => n8469, B2 => 
                           n9755, ZN => n3475);
   U1894 : OAI22_X1 port map( A1 => n9238, A2 => n9746, B1 => n8470, B2 => 
                           n9755, ZN => n3459);
   U1895 : OAI22_X1 port map( A1 => n9331, A2 => n9736, B1 => n8510, B2 => 
                           n9737, ZN => n3954);
   U1896 : OAI22_X1 port map( A1 => n9328, A2 => n9735, B1 => n8511, B2 => 
                           n9737, ZN => n3938);
   U1897 : OAI22_X1 port map( A1 => n9325, A2 => n9736, B1 => n8512, B2 => 
                           n9737, ZN => n3922);
   U1898 : OAI22_X1 port map( A1 => n9322, A2 => n9735, B1 => n8513, B2 => 
                           n9737, ZN => n3906);
   U1899 : OAI22_X1 port map( A1 => n9319, A2 => n9736, B1 => n8514, B2 => 
                           n9738, ZN => n3890);
   U1900 : OAI22_X1 port map( A1 => n9316, A2 => n9735, B1 => n8515, B2 => 
                           n9738, ZN => n3874);
   U1901 : OAI22_X1 port map( A1 => n9313, A2 => n9736, B1 => n8516, B2 => 
                           n9738, ZN => n3858);
   U1902 : OAI22_X1 port map( A1 => n9310, A2 => n9735, B1 => n8517, B2 => 
                           n9738, ZN => n3842);
   U1903 : OAI22_X1 port map( A1 => n9307, A2 => n9736, B1 => n8518, B2 => 
                           n9739, ZN => n3826);
   U1904 : OAI22_X1 port map( A1 => n9304, A2 => n9736, B1 => n8519, B2 => 
                           n9739, ZN => n3810);
   U1905 : OAI22_X1 port map( A1 => n9301, A2 => n9736, B1 => n8520, B2 => 
                           n9739, ZN => n3794);
   U1906 : OAI22_X1 port map( A1 => n9298, A2 => n9736, B1 => n8521, B2 => 
                           n9739, ZN => n3778);
   U1907 : OAI22_X1 port map( A1 => n9295, A2 => n9736, B1 => n8522, B2 => 
                           n9740, ZN => n3762);
   U1908 : OAI22_X1 port map( A1 => n9292, A2 => n9736, B1 => n8523, B2 => 
                           n9740, ZN => n3746);
   U1909 : OAI22_X1 port map( A1 => n9289, A2 => n9736, B1 => n8524, B2 => 
                           n9740, ZN => n3730);
   U1910 : OAI22_X1 port map( A1 => n9286, A2 => n9736, B1 => n8525, B2 => 
                           n9740, ZN => n3714);
   U1911 : OAI22_X1 port map( A1 => n9283, A2 => n9736, B1 => n8526, B2 => 
                           n9741, ZN => n3698);
   U1912 : OAI22_X1 port map( A1 => n9280, A2 => n9736, B1 => n8527, B2 => 
                           n9741, ZN => n3682);
   U1913 : OAI22_X1 port map( A1 => n9277, A2 => n9736, B1 => n8528, B2 => 
                           n9741, ZN => n3666);
   U1914 : OAI22_X1 port map( A1 => n9274, A2 => n9736, B1 => n8529, B2 => 
                           n9741, ZN => n3650);
   U1915 : OAI22_X1 port map( A1 => n9271, A2 => n9735, B1 => n8530, B2 => 
                           n9742, ZN => n3634);
   U1916 : OAI22_X1 port map( A1 => n9268, A2 => n9735, B1 => n8531, B2 => 
                           n9742, ZN => n3618);
   U1917 : OAI22_X1 port map( A1 => n9265, A2 => n9735, B1 => n8532, B2 => 
                           n9742, ZN => n3602);
   U1918 : OAI22_X1 port map( A1 => n9262, A2 => n9735, B1 => n8533, B2 => 
                           n9742, ZN => n3586);
   U1919 : OAI22_X1 port map( A1 => n9259, A2 => n9735, B1 => n8534, B2 => 
                           n9743, ZN => n3570);
   U1920 : OAI22_X1 port map( A1 => n9256, A2 => n9735, B1 => n8535, B2 => 
                           n9743, ZN => n3554);
   U1921 : OAI22_X1 port map( A1 => n9253, A2 => n9735, B1 => n8536, B2 => 
                           n9743, ZN => n3538);
   U1922 : OAI22_X1 port map( A1 => n9250, A2 => n9735, B1 => n8537, B2 => 
                           n9743, ZN => n3522);
   U1923 : OAI22_X1 port map( A1 => n9247, A2 => n9735, B1 => n8538, B2 => 
                           n9744, ZN => n3506);
   U1924 : OAI22_X1 port map( A1 => n9244, A2 => n9735, B1 => n8539, B2 => 
                           n9744, ZN => n3490);
   U1925 : OAI22_X1 port map( A1 => n9241, A2 => n9735, B1 => n8540, B2 => 
                           n9744, ZN => n3474);
   U1926 : OAI22_X1 port map( A1 => n9238, A2 => n9735, B1 => n8541, B2 => 
                           n9744, ZN => n3458);
   U1927 : OAI22_X1 port map( A1 => n9329, A2 => n9725, B1 => n8599, B2 => 
                           n9726, ZN => n3936);
   U1928 : OAI22_X1 port map( A1 => n9326, A2 => n9724, B1 => n8600, B2 => 
                           n9726, ZN => n3920);
   U1929 : OAI22_X1 port map( A1 => n9323, A2 => n9725, B1 => n8601, B2 => 
                           n9726, ZN => n3904);
   U1930 : OAI22_X1 port map( A1 => n9320, A2 => n9724, B1 => n8602, B2 => 
                           n9727, ZN => n3888);
   U1931 : OAI22_X1 port map( A1 => n9317, A2 => n9725, B1 => n8603, B2 => 
                           n9727, ZN => n3872);
   U1932 : OAI22_X1 port map( A1 => n9314, A2 => n9724, B1 => n8604, B2 => 
                           n9727, ZN => n3856);
   U1933 : OAI22_X1 port map( A1 => n9311, A2 => n9725, B1 => n8605, B2 => 
                           n9727, ZN => n3840);
   U1934 : OAI22_X1 port map( A1 => n9308, A2 => n9725, B1 => n8606, B2 => 
                           n9728, ZN => n3824);
   U1935 : OAI22_X1 port map( A1 => n9305, A2 => n9725, B1 => n8607, B2 => 
                           n9728, ZN => n3808);
   U1936 : OAI22_X1 port map( A1 => n9302, A2 => n9725, B1 => n8608, B2 => 
                           n9728, ZN => n3792);
   U1937 : OAI22_X1 port map( A1 => n9299, A2 => n9725, B1 => n8609, B2 => 
                           n9728, ZN => n3776);
   U1938 : OAI22_X1 port map( A1 => n9296, A2 => n9725, B1 => n8610, B2 => 
                           n9729, ZN => n3760);
   U1939 : OAI22_X1 port map( A1 => n9293, A2 => n9725, B1 => n8611, B2 => 
                           n9729, ZN => n3744);
   U1940 : OAI22_X1 port map( A1 => n9290, A2 => n9725, B1 => n8612, B2 => 
                           n9729, ZN => n3728);
   U1941 : OAI22_X1 port map( A1 => n9287, A2 => n9725, B1 => n8613, B2 => 
                           n9729, ZN => n3712);
   U1942 : OAI22_X1 port map( A1 => n9284, A2 => n9725, B1 => n8614, B2 => 
                           n9730, ZN => n3696);
   U1943 : OAI22_X1 port map( A1 => n9281, A2 => n9725, B1 => n8615, B2 => 
                           n9730, ZN => n3680);
   U1944 : OAI22_X1 port map( A1 => n9278, A2 => n9725, B1 => n8616, B2 => 
                           n9730, ZN => n3664);
   U1945 : OAI22_X1 port map( A1 => n9275, A2 => n9725, B1 => n8617, B2 => 
                           n9730, ZN => n3648);
   U1946 : OAI22_X1 port map( A1 => n9272, A2 => n9724, B1 => n8618, B2 => 
                           n9731, ZN => n3632);
   U1947 : OAI22_X1 port map( A1 => n9269, A2 => n9724, B1 => n8619, B2 => 
                           n9731, ZN => n3616);
   U1948 : OAI22_X1 port map( A1 => n9266, A2 => n9724, B1 => n8620, B2 => 
                           n9731, ZN => n3600);
   U1949 : OAI22_X1 port map( A1 => n9263, A2 => n9724, B1 => n8621, B2 => 
                           n9731, ZN => n3584);
   U1950 : OAI22_X1 port map( A1 => n9260, A2 => n9724, B1 => n8622, B2 => 
                           n9732, ZN => n3568);
   U1951 : OAI22_X1 port map( A1 => n9257, A2 => n9724, B1 => n8623, B2 => 
                           n9732, ZN => n3552);
   U1952 : OAI22_X1 port map( A1 => n9254, A2 => n9724, B1 => n8624, B2 => 
                           n9732, ZN => n3536);
   U1953 : OAI22_X1 port map( A1 => n9251, A2 => n9724, B1 => n8625, B2 => 
                           n9732, ZN => n3520);
   U1954 : OAI22_X1 port map( A1 => n9248, A2 => n9724, B1 => n8626, B2 => 
                           n9733, ZN => n3504);
   U1955 : OAI22_X1 port map( A1 => n9245, A2 => n9724, B1 => n8627, B2 => 
                           n9733, ZN => n3488);
   U1956 : OAI22_X1 port map( A1 => n9242, A2 => n9724, B1 => n8628, B2 => 
                           n9733, ZN => n3472);
   U1957 : OAI22_X1 port map( A1 => n9239, A2 => n9724, B1 => n8629, B2 => 
                           n9733, ZN => n3456);
   U1958 : OAI22_X1 port map( A1 => n9332, A2 => n9625, B1 => n8742, B2 => 
                           n9634, ZN => n3262);
   U1959 : OAI22_X1 port map( A1 => n9329, A2 => n9625, B1 => n8743, B2 => 
                           n9634, ZN => n3263);
   U1960 : OAI22_X1 port map( A1 => n9326, A2 => n9625, B1 => n8744, B2 => 
                           n9634, ZN => n3264);
   U1961 : OAI22_X1 port map( A1 => n9323, A2 => n9625, B1 => n8745, B2 => 
                           n9634, ZN => n3265);
   U1962 : OAI22_X1 port map( A1 => n9320, A2 => n9625, B1 => n8746, B2 => 
                           n9633, ZN => n3266);
   U1963 : OAI22_X1 port map( A1 => n9317, A2 => n9625, B1 => n8747, B2 => 
                           n9633, ZN => n3267);
   U1964 : OAI22_X1 port map( A1 => n9314, A2 => n9625, B1 => n8748, B2 => 
                           n9633, ZN => n3268);
   U1965 : OAI22_X1 port map( A1 => n9311, A2 => n9625, B1 => n8749, B2 => 
                           n9633, ZN => n3269);
   U1966 : OAI22_X1 port map( A1 => n9308, A2 => n9625, B1 => n8750, B2 => 
                           n9632, ZN => n3270);
   U1967 : OAI22_X1 port map( A1 => n9305, A2 => n9625, B1 => n8751, B2 => 
                           n9632, ZN => n3271);
   U1968 : OAI22_X1 port map( A1 => n9302, A2 => n9625, B1 => n8752, B2 => 
                           n9632, ZN => n3272);
   U1969 : OAI22_X1 port map( A1 => n9299, A2 => n9625, B1 => n8753, B2 => 
                           n9632, ZN => n3273);
   U1970 : OAI22_X1 port map( A1 => n9296, A2 => n9626, B1 => n8754, B2 => 
                           n9631, ZN => n3274);
   U1971 : OAI22_X1 port map( A1 => n9293, A2 => n9626, B1 => n8755, B2 => 
                           n9631, ZN => n3275);
   U1972 : OAI22_X1 port map( A1 => n9290, A2 => n9626, B1 => n8756, B2 => 
                           n9631, ZN => n3276);
   U1973 : OAI22_X1 port map( A1 => n9287, A2 => n9626, B1 => n8757, B2 => 
                           n9631, ZN => n3277);
   U1974 : OAI22_X1 port map( A1 => n9284, A2 => n9626, B1 => n8758, B2 => 
                           n9630, ZN => n3278);
   U1975 : OAI22_X1 port map( A1 => n9281, A2 => n9626, B1 => n8759, B2 => 
                           n9630, ZN => n3279);
   U1976 : OAI22_X1 port map( A1 => n9278, A2 => n9626, B1 => n8760, B2 => 
                           n9630, ZN => n3280);
   U1977 : OAI22_X1 port map( A1 => n9275, A2 => n9626, B1 => n8761, B2 => 
                           n9630, ZN => n3281);
   U1978 : OAI22_X1 port map( A1 => n9272, A2 => n9626, B1 => n8762, B2 => 
                           n9629, ZN => n3282);
   U1979 : OAI22_X1 port map( A1 => n9269, A2 => n9626, B1 => n8763, B2 => 
                           n9629, ZN => n3283);
   U1980 : OAI22_X1 port map( A1 => n9266, A2 => n9626, B1 => n8764, B2 => 
                           n9629, ZN => n3284);
   U1981 : OAI22_X1 port map( A1 => n9263, A2 => n9626, B1 => n8765, B2 => 
                           n9629, ZN => n3285);
   U1982 : OAI22_X1 port map( A1 => n9260, A2 => n9625, B1 => n8766, B2 => 
                           n9628, ZN => n3286);
   U1983 : OAI22_X1 port map( A1 => n9257, A2 => n9626, B1 => n8767, B2 => 
                           n9628, ZN => n3287);
   U1984 : OAI22_X1 port map( A1 => n9254, A2 => n9625, B1 => n8768, B2 => 
                           n9628, ZN => n3288);
   U1985 : OAI22_X1 port map( A1 => n9251, A2 => n9626, B1 => n8769, B2 => 
                           n9628, ZN => n3289);
   U1986 : OAI22_X1 port map( A1 => n9248, A2 => n9625, B1 => n8770, B2 => 
                           n9627, ZN => n3290);
   U1987 : OAI22_X1 port map( A1 => n9245, A2 => n9626, B1 => n8771, B2 => 
                           n9627, ZN => n3291);
   U1988 : OAI22_X1 port map( A1 => n9242, A2 => n9625, B1 => n8772, B2 => 
                           n9627, ZN => n3292);
   U1989 : OAI22_X1 port map( A1 => n9239, A2 => n9626, B1 => n8773, B2 => 
                           n9627, ZN => n3293);
   U1990 : OAI22_X1 port map( A1 => n9332, A2 => n9692, B1 => n8830, B2 => 
                           n9693, ZN => n3946);
   U1991 : OAI22_X1 port map( A1 => n9329, A2 => n9691, B1 => n8831, B2 => 
                           n9693, ZN => n3930);
   U1992 : OAI22_X1 port map( A1 => n9326, A2 => n9692, B1 => n8832, B2 => 
                           n9693, ZN => n3914);
   U1993 : OAI22_X1 port map( A1 => n9323, A2 => n9691, B1 => n8833, B2 => 
                           n9693, ZN => n3898);
   U1994 : OAI22_X1 port map( A1 => n9320, A2 => n9692, B1 => n8834, B2 => 
                           n9694, ZN => n3882);
   U1995 : OAI22_X1 port map( A1 => n9317, A2 => n9691, B1 => n8835, B2 => 
                           n9694, ZN => n3866);
   U1996 : OAI22_X1 port map( A1 => n9314, A2 => n9692, B1 => n8836, B2 => 
                           n9694, ZN => n3850);
   U1997 : OAI22_X1 port map( A1 => n9311, A2 => n9691, B1 => n8837, B2 => 
                           n9694, ZN => n3834);
   U1998 : OAI22_X1 port map( A1 => n9308, A2 => n9692, B1 => n8838, B2 => 
                           n9695, ZN => n3818);
   U1999 : OAI22_X1 port map( A1 => n9305, A2 => n9692, B1 => n8839, B2 => 
                           n9695, ZN => n3802);
   U2000 : OAI22_X1 port map( A1 => n9302, A2 => n9692, B1 => n8840, B2 => 
                           n9695, ZN => n3786);
   U2001 : OAI22_X1 port map( A1 => n9299, A2 => n9692, B1 => n8841, B2 => 
                           n9695, ZN => n3770);
   U2002 : OAI22_X1 port map( A1 => n9296, A2 => n9692, B1 => n8842, B2 => 
                           n9696, ZN => n3754);
   U2003 : OAI22_X1 port map( A1 => n9293, A2 => n9692, B1 => n8843, B2 => 
                           n9696, ZN => n3738);
   U2004 : OAI22_X1 port map( A1 => n9290, A2 => n9692, B1 => n8844, B2 => 
                           n9696, ZN => n3722);
   U2005 : OAI22_X1 port map( A1 => n9287, A2 => n9692, B1 => n8845, B2 => 
                           n9696, ZN => n3706);
   U2006 : OAI22_X1 port map( A1 => n9284, A2 => n9692, B1 => n8846, B2 => 
                           n9697, ZN => n3690);
   U2007 : OAI22_X1 port map( A1 => n9281, A2 => n9692, B1 => n8847, B2 => 
                           n9697, ZN => n3674);
   U2008 : OAI22_X1 port map( A1 => n9278, A2 => n9692, B1 => n8848, B2 => 
                           n9697, ZN => n3658);
   U2009 : OAI22_X1 port map( A1 => n9275, A2 => n9692, B1 => n8849, B2 => 
                           n9697, ZN => n3642);
   U2010 : OAI22_X1 port map( A1 => n9272, A2 => n9691, B1 => n8850, B2 => 
                           n9698, ZN => n3626);
   U2011 : OAI22_X1 port map( A1 => n9269, A2 => n9691, B1 => n8851, B2 => 
                           n9698, ZN => n3610);
   U2012 : OAI22_X1 port map( A1 => n9266, A2 => n9691, B1 => n8852, B2 => 
                           n9698, ZN => n3594);
   U2013 : OAI22_X1 port map( A1 => n9263, A2 => n9691, B1 => n8853, B2 => 
                           n9698, ZN => n3578);
   U2014 : OAI22_X1 port map( A1 => n9260, A2 => n9691, B1 => n8854, B2 => 
                           n9699, ZN => n3562);
   U2015 : OAI22_X1 port map( A1 => n9257, A2 => n9691, B1 => n8855, B2 => 
                           n9699, ZN => n3546);
   U2016 : OAI22_X1 port map( A1 => n9254, A2 => n9691, B1 => n8856, B2 => 
                           n9699, ZN => n3530);
   U2017 : OAI22_X1 port map( A1 => n9251, A2 => n9691, B1 => n8857, B2 => 
                           n9699, ZN => n3514);
   U2018 : OAI22_X1 port map( A1 => n9248, A2 => n9691, B1 => n8858, B2 => 
                           n9700, ZN => n3498);
   U2019 : OAI22_X1 port map( A1 => n9245, A2 => n9691, B1 => n8859, B2 => 
                           n9700, ZN => n3482);
   U2020 : OAI22_X1 port map( A1 => n9242, A2 => n9691, B1 => n8860, B2 => 
                           n9700, ZN => n3466);
   U2021 : OAI22_X1 port map( A1 => n9239, A2 => n9691, B1 => n8861, B2 => 
                           n9700, ZN => n3450);
   U2022 : OAI22_X1 port map( A1 => n9332, A2 => n9681, B1 => n8918, B2 => 
                           n9682, ZN => n3944);
   U2023 : OAI22_X1 port map( A1 => n9329, A2 => n9680, B1 => n8919, B2 => 
                           n9682, ZN => n3928);
   U2024 : OAI22_X1 port map( A1 => n9326, A2 => n9681, B1 => n8920, B2 => 
                           n9682, ZN => n3912);
   U2025 : OAI22_X1 port map( A1 => n9323, A2 => n9680, B1 => n8921, B2 => 
                           n9682, ZN => n3896);
   U2026 : OAI22_X1 port map( A1 => n9320, A2 => n9681, B1 => n8922, B2 => 
                           n9683, ZN => n3880);
   U2027 : OAI22_X1 port map( A1 => n9317, A2 => n9680, B1 => n8923, B2 => 
                           n9683, ZN => n3864);
   U2028 : OAI22_X1 port map( A1 => n9314, A2 => n9681, B1 => n8924, B2 => 
                           n9683, ZN => n3848);
   U2029 : OAI22_X1 port map( A1 => n9311, A2 => n9680, B1 => n8925, B2 => 
                           n9683, ZN => n3832);
   U2030 : OAI22_X1 port map( A1 => n9308, A2 => n9681, B1 => n8926, B2 => 
                           n9684, ZN => n3816);
   U2031 : OAI22_X1 port map( A1 => n9305, A2 => n9681, B1 => n8927, B2 => 
                           n9684, ZN => n3800);
   U2032 : OAI22_X1 port map( A1 => n9302, A2 => n9681, B1 => n8928, B2 => 
                           n9684, ZN => n3784);
   U2033 : OAI22_X1 port map( A1 => n9299, A2 => n9681, B1 => n8929, B2 => 
                           n9684, ZN => n3768);
   U2034 : OAI22_X1 port map( A1 => n9296, A2 => n9681, B1 => n8930, B2 => 
                           n9685, ZN => n3752);
   U2035 : OAI22_X1 port map( A1 => n9293, A2 => n9681, B1 => n8931, B2 => 
                           n9685, ZN => n3736);
   U2036 : OAI22_X1 port map( A1 => n9290, A2 => n9681, B1 => n8932, B2 => 
                           n9685, ZN => n3720);
   U2037 : OAI22_X1 port map( A1 => n9287, A2 => n9681, B1 => n8933, B2 => 
                           n9685, ZN => n3704);
   U2038 : OAI22_X1 port map( A1 => n9284, A2 => n9681, B1 => n8934, B2 => 
                           n9686, ZN => n3688);
   U2039 : OAI22_X1 port map( A1 => n9281, A2 => n9681, B1 => n8935, B2 => 
                           n9686, ZN => n3672);
   U2040 : OAI22_X1 port map( A1 => n9278, A2 => n9681, B1 => n8936, B2 => 
                           n9686, ZN => n3656);
   U2041 : OAI22_X1 port map( A1 => n9275, A2 => n9681, B1 => n8937, B2 => 
                           n9686, ZN => n3640);
   U2042 : OAI22_X1 port map( A1 => n9272, A2 => n9680, B1 => n8938, B2 => 
                           n9687, ZN => n3624);
   U2043 : OAI22_X1 port map( A1 => n9269, A2 => n9680, B1 => n8939, B2 => 
                           n9687, ZN => n3608);
   U2044 : OAI22_X1 port map( A1 => n9266, A2 => n9680, B1 => n8940, B2 => 
                           n9687, ZN => n3592);
   U2045 : OAI22_X1 port map( A1 => n9263, A2 => n9680, B1 => n8941, B2 => 
                           n9687, ZN => n3576);
   U2046 : OAI22_X1 port map( A1 => n9260, A2 => n9680, B1 => n8942, B2 => 
                           n9688, ZN => n3560);
   U2047 : OAI22_X1 port map( A1 => n9257, A2 => n9680, B1 => n8943, B2 => 
                           n9688, ZN => n3544);
   U2048 : OAI22_X1 port map( A1 => n9254, A2 => n9680, B1 => n8944, B2 => 
                           n9688, ZN => n3528);
   U2049 : OAI22_X1 port map( A1 => n9251, A2 => n9680, B1 => n8945, B2 => 
                           n9688, ZN => n3512);
   U2050 : OAI22_X1 port map( A1 => n9248, A2 => n9680, B1 => n8946, B2 => 
                           n9689, ZN => n3496);
   U2051 : OAI22_X1 port map( A1 => n9245, A2 => n9680, B1 => n8947, B2 => 
                           n9689, ZN => n3480);
   U2052 : OAI22_X1 port map( A1 => n9242, A2 => n9680, B1 => n8948, B2 => 
                           n9689, ZN => n3464);
   U2053 : OAI22_X1 port map( A1 => n9239, A2 => n9680, B1 => n8949, B2 => 
                           n9689, ZN => n3448);
   U2054 : OAI22_X1 port map( A1 => n9875, A2 => n9331, B1 => n2349, B2 => 
                           n9867, ZN => n9174);
   U2055 : OAI22_X1 port map( A1 => n9875, A2 => n9328, B1 => n2341, B2 => 
                           n9867, ZN => n9175);
   U2056 : OAI22_X1 port map( A1 => n9874, A2 => n9325, B1 => n2333, B2 => 
                           n9867, ZN => n9176);
   U2057 : OAI22_X1 port map( A1 => n9874, A2 => n9322, B1 => n2325, B2 => 
                           n9867, ZN => n9177);
   U2058 : OAI22_X1 port map( A1 => n9874, A2 => n9319, B1 => n2317, B2 => 
                           n9867, ZN => n9178);
   U2059 : OAI22_X1 port map( A1 => n9874, A2 => n9316, B1 => n2309, B2 => 
                           n9867, ZN => n9179);
   U2060 : OAI22_X1 port map( A1 => n9874, A2 => n9313, B1 => n2301, B2 => 
                           n9867, ZN => n9180);
   U2061 : OAI22_X1 port map( A1 => n9873, A2 => n9310, B1 => n2293, B2 => 
                           n9867, ZN => n9181);
   U2062 : OAI22_X1 port map( A1 => n9873, A2 => n9307, B1 => n2285, B2 => 
                           n9867, ZN => n9182);
   U2063 : OAI22_X1 port map( A1 => n9873, A2 => n9304, B1 => n2277, B2 => 
                           n9867, ZN => n9183);
   U2064 : OAI22_X1 port map( A1 => n9873, A2 => n9301, B1 => n2269, B2 => 
                           n9867, ZN => n9184);
   U2065 : OAI22_X1 port map( A1 => n9873, A2 => n9298, B1 => n2261, B2 => 
                           n9867, ZN => n9185);
   U2066 : OAI22_X1 port map( A1 => n9872, A2 => n9295, B1 => n2253, B2 => 
                           n9868, ZN => n9186);
   U2067 : OAI22_X1 port map( A1 => n9872, A2 => n9292, B1 => n2245, B2 => 
                           n9868, ZN => n9187);
   U2068 : OAI22_X1 port map( A1 => n9872, A2 => n9289, B1 => n2237, B2 => 
                           n9868, ZN => n9188);
   U2069 : OAI22_X1 port map( A1 => n9872, A2 => n9286, B1 => n2229, B2 => 
                           n9868, ZN => n9189);
   U2070 : OAI22_X1 port map( A1 => n9872, A2 => n9283, B1 => n2221, B2 => 
                           n9868, ZN => n9190);
   U2071 : OAI22_X1 port map( A1 => n9871, A2 => n9280, B1 => n2213, B2 => 
                           n9868, ZN => n9191);
   U2072 : OAI22_X1 port map( A1 => n9871, A2 => n9277, B1 => n2205, B2 => 
                           n9868, ZN => n9192);
   U2073 : OAI22_X1 port map( A1 => n9871, A2 => n9274, B1 => n2197, B2 => 
                           n9868, ZN => n9193);
   U2074 : OAI22_X1 port map( A1 => n9871, A2 => n9271, B1 => n2189, B2 => 
                           n9868, ZN => n9194);
   U2075 : OAI22_X1 port map( A1 => n9871, A2 => n9268, B1 => n2181, B2 => 
                           n9868, ZN => n9195);
   U2076 : OAI22_X1 port map( A1 => n9870, A2 => n9265, B1 => n2173, B2 => 
                           n9868, ZN => n9196);
   U2077 : OAI22_X1 port map( A1 => n9870, A2 => n9262, B1 => n2165, B2 => 
                           n9868, ZN => n9197);
   U2078 : OAI22_X1 port map( A1 => n9312, A2 => n9548, B1 => n8246, B2 => 
                           n9556, ZN => n3045);
   U2079 : OAI22_X1 port map( A1 => n9309, A2 => n9548, B1 => n8247, B2 => 
                           n9555, ZN => n3046);
   U2080 : OAI22_X1 port map( A1 => n9306, A2 => n9548, B1 => n8248, B2 => 
                           n9555, ZN => n3047);
   U2081 : OAI22_X1 port map( A1 => n9303, A2 => n9548, B1 => n8249, B2 => 
                           n9555, ZN => n3048);
   U2082 : OAI22_X1 port map( A1 => n9300, A2 => n9548, B1 => n8250, B2 => 
                           n9555, ZN => n3049);
   U2083 : OAI22_X1 port map( A1 => n9297, A2 => n9549, B1 => n8251, B2 => 
                           n9554, ZN => n3050);
   U2084 : OAI22_X1 port map( A1 => n9294, A2 => n9549, B1 => n8252, B2 => 
                           n9554, ZN => n3051);
   U2085 : OAI22_X1 port map( A1 => n9291, A2 => n9549, B1 => n8253, B2 => 
                           n9554, ZN => n3052);
   U2086 : OAI22_X1 port map( A1 => n9288, A2 => n9549, B1 => n8254, B2 => 
                           n9554, ZN => n3053);
   U2087 : OAI22_X1 port map( A1 => n9285, A2 => n9549, B1 => n8255, B2 => 
                           n9553, ZN => n3054);
   U2088 : OAI22_X1 port map( A1 => n9282, A2 => n9549, B1 => n8256, B2 => 
                           n9553, ZN => n3055);
   U2089 : OAI22_X1 port map( A1 => n9279, A2 => n9549, B1 => n8257, B2 => 
                           n9553, ZN => n3056);
   U2090 : OAI22_X1 port map( A1 => n9276, A2 => n9549, B1 => n8258, B2 => 
                           n9553, ZN => n3057);
   U2091 : OAI22_X1 port map( A1 => n9273, A2 => n9549, B1 => n8259, B2 => 
                           n9552, ZN => n3058);
   U2092 : OAI22_X1 port map( A1 => n9270, A2 => n9549, B1 => n8260, B2 => 
                           n9552, ZN => n3059);
   U2093 : OAI22_X1 port map( A1 => n9267, A2 => n9549, B1 => n8261, B2 => 
                           n9552, ZN => n3060);
   U2094 : OAI22_X1 port map( A1 => n9264, A2 => n9549, B1 => n8262, B2 => 
                           n9552, ZN => n3061);
   U2095 : OAI22_X1 port map( A1 => n9260, A2 => n9636, B1 => n8311, B2 => 
                           n9639, ZN => n3318);
   U2096 : OAI22_X1 port map( A1 => n9257, A2 => n9637, B1 => n8312, B2 => 
                           n9639, ZN => n3319);
   U2097 : OAI22_X1 port map( A1 => n9254, A2 => n9636, B1 => n8313, B2 => 
                           n9639, ZN => n3320);
   U2098 : OAI22_X1 port map( A1 => n9251, A2 => n9637, B1 => n8314, B2 => 
                           n9639, ZN => n3321);
   U2099 : OAI22_X1 port map( A1 => n9248, A2 => n9636, B1 => n8315, B2 => 
                           n9638, ZN => n3322);
   U2100 : OAI22_X1 port map( A1 => n9245, A2 => n9637, B1 => n8316, B2 => 
                           n9638, ZN => n3323);
   U2101 : OAI22_X1 port map( A1 => n9242, A2 => n9636, B1 => n8317, B2 => 
                           n9638, ZN => n3324);
   U2102 : OAI22_X1 port map( A1 => n9239, A2 => n9637, B1 => n8318, B2 => 
                           n9638, ZN => n3325);
   U2103 : OAI22_X1 port map( A1 => n9261, A2 => n9549, B1 => n8327, B2 => 
                           n9551, ZN => n3062);
   U2104 : OAI22_X1 port map( A1 => n9258, A2 => n9548, B1 => n8328, B2 => 
                           n9551, ZN => n3063);
   U2105 : OAI22_X1 port map( A1 => n9255, A2 => n9549, B1 => n8329, B2 => 
                           n9551, ZN => n3064);
   U2106 : OAI22_X1 port map( A1 => n9252, A2 => n9548, B1 => n8330, B2 => 
                           n9551, ZN => n3065);
   U2107 : OAI22_X1 port map( A1 => n9249, A2 => n9549, B1 => n8331, B2 => 
                           n9550, ZN => n3066);
   U2108 : OAI22_X1 port map( A1 => n9246, A2 => n9548, B1 => n8332, B2 => 
                           n9550, ZN => n3067);
   U2109 : OAI22_X1 port map( A1 => n9243, A2 => n9549, B1 => n8333, B2 => 
                           n9550, ZN => n3068);
   U2110 : OAI22_X1 port map( A1 => n9240, A2 => n9548, B1 => n8334, B2 => 
                           n9550, ZN => n3069);
   U2111 : OAI22_X1 port map( A1 => n9331, A2 => n9769, B1 => n8375, B2 => 
                           n9770, ZN => n3957);
   U2112 : OAI22_X1 port map( A1 => n9328, A2 => n9768, B1 => n8376, B2 => 
                           n9770, ZN => n3941);
   U2113 : OAI22_X1 port map( A1 => n9325, A2 => n9769, B1 => n8377, B2 => 
                           n9770, ZN => n3925);
   U2114 : OAI22_X1 port map( A1 => n9322, A2 => n9768, B1 => n8378, B2 => 
                           n9770, ZN => n3909);
   U2115 : OAI22_X1 port map( A1 => n9319, A2 => n9769, B1 => n8379, B2 => 
                           n9771, ZN => n3893);
   U2116 : OAI22_X1 port map( A1 => n9316, A2 => n9768, B1 => n8380, B2 => 
                           n9771, ZN => n3877);
   U2117 : OAI22_X1 port map( A1 => n9313, A2 => n9769, B1 => n8381, B2 => 
                           n9771, ZN => n3861);
   U2118 : OAI22_X1 port map( A1 => n9310, A2 => n9768, B1 => n8382, B2 => 
                           n9771, ZN => n3845);
   U2119 : OAI22_X1 port map( A1 => n9307, A2 => n9769, B1 => n8383, B2 => 
                           n9772, ZN => n3829);
   U2120 : OAI22_X1 port map( A1 => n9304, A2 => n9769, B1 => n8384, B2 => 
                           n9772, ZN => n3813);
   U2121 : OAI22_X1 port map( A1 => n9301, A2 => n9769, B1 => n8385, B2 => 
                           n9772, ZN => n3797);
   U2122 : OAI22_X1 port map( A1 => n9298, A2 => n9769, B1 => n8386, B2 => 
                           n9772, ZN => n3781);
   U2123 : OAI22_X1 port map( A1 => n9295, A2 => n9769, B1 => n8387, B2 => 
                           n9773, ZN => n3765);
   U2124 : OAI22_X1 port map( A1 => n9292, A2 => n9769, B1 => n8388, B2 => 
                           n9773, ZN => n3749);
   U2125 : OAI22_X1 port map( A1 => n9289, A2 => n9769, B1 => n8389, B2 => 
                           n9773, ZN => n3733);
   U2126 : OAI22_X1 port map( A1 => n9286, A2 => n9769, B1 => n8390, B2 => 
                           n9773, ZN => n3717);
   U2127 : OAI22_X1 port map( A1 => n9283, A2 => n9769, B1 => n8391, B2 => 
                           n9774, ZN => n3701);
   U2128 : OAI22_X1 port map( A1 => n9280, A2 => n9769, B1 => n8392, B2 => 
                           n9774, ZN => n3685);
   U2129 : OAI22_X1 port map( A1 => n9277, A2 => n9769, B1 => n8393, B2 => 
                           n9774, ZN => n3669);
   U2130 : OAI22_X1 port map( A1 => n9274, A2 => n9769, B1 => n8394, B2 => 
                           n9774, ZN => n3653);
   U2131 : OAI22_X1 port map( A1 => n9271, A2 => n9768, B1 => n8395, B2 => 
                           n9775, ZN => n3637);
   U2132 : OAI22_X1 port map( A1 => n9268, A2 => n9768, B1 => n8396, B2 => 
                           n9775, ZN => n3621);
   U2133 : OAI22_X1 port map( A1 => n9265, A2 => n9768, B1 => n8397, B2 => 
                           n9775, ZN => n3605);
   U2134 : OAI22_X1 port map( A1 => n9262, A2 => n9768, B1 => n8398, B2 => 
                           n9775, ZN => n3589);
   U2135 : OAI22_X1 port map( A1 => n9259, A2 => n9768, B1 => n8399, B2 => 
                           n9776, ZN => n3573);
   U2136 : OAI22_X1 port map( A1 => n9256, A2 => n9768, B1 => n8400, B2 => 
                           n9776, ZN => n3557);
   U2137 : OAI22_X1 port map( A1 => n9253, A2 => n9768, B1 => n8401, B2 => 
                           n9776, ZN => n3541);
   U2138 : OAI22_X1 port map( A1 => n9250, A2 => n9768, B1 => n8402, B2 => 
                           n9776, ZN => n3525);
   U2139 : OAI22_X1 port map( A1 => n9247, A2 => n9768, B1 => n8403, B2 => 
                           n9777, ZN => n3509);
   U2140 : OAI22_X1 port map( A1 => n9244, A2 => n9768, B1 => n8404, B2 => 
                           n9777, ZN => n3493);
   U2141 : OAI22_X1 port map( A1 => n9241, A2 => n9768, B1 => n8405, B2 => 
                           n9777, ZN => n3477);
   U2142 : OAI22_X1 port map( A1 => n9238, A2 => n9768, B1 => n8406, B2 => 
                           n9777, ZN => n3461);
   U2143 : OAI22_X1 port map( A1 => n9333, A2 => n9548, B1 => n8471, B2 => 
                           n9557, ZN => n3038);
   U2144 : OAI22_X1 port map( A1 => n9330, A2 => n9548, B1 => n8472, B2 => 
                           n9557, ZN => n3039);
   U2145 : OAI22_X1 port map( A1 => n9327, A2 => n9548, B1 => n8473, B2 => 
                           n9557, ZN => n3040);
   U2146 : OAI22_X1 port map( A1 => n9324, A2 => n9548, B1 => n8474, B2 => 
                           n9557, ZN => n3041);
   U2147 : OAI22_X1 port map( A1 => n9321, A2 => n9548, B1 => n8475, B2 => 
                           n9556, ZN => n3042);
   U2148 : OAI22_X1 port map( A1 => n9318, A2 => n9548, B1 => n8476, B2 => 
                           n9556, ZN => n3043);
   U2149 : OAI22_X1 port map( A1 => n9315, A2 => n9548, B1 => n8477, B2 => 
                           n9556, ZN => n3044);
   U2150 : OAI22_X1 port map( A1 => n9333, A2 => n9559, B1 => n8478, B2 => 
                           n9568, ZN => n3070);
   U2151 : OAI22_X1 port map( A1 => n9330, A2 => n9559, B1 => n8479, B2 => 
                           n9568, ZN => n3071);
   U2152 : OAI22_X1 port map( A1 => n9327, A2 => n9559, B1 => n8480, B2 => 
                           n9568, ZN => n3072);
   U2153 : OAI22_X1 port map( A1 => n9324, A2 => n9559, B1 => n8481, B2 => 
                           n9568, ZN => n3073);
   U2154 : OAI22_X1 port map( A1 => n9321, A2 => n9559, B1 => n8482, B2 => 
                           n9567, ZN => n3074);
   U2155 : OAI22_X1 port map( A1 => n9318, A2 => n9559, B1 => n8483, B2 => 
                           n9567, ZN => n3075);
   U2156 : OAI22_X1 port map( A1 => n9315, A2 => n9559, B1 => n8484, B2 => 
                           n9567, ZN => n3076);
   U2157 : OAI22_X1 port map( A1 => n9312, A2 => n9559, B1 => n8485, B2 => 
                           n9567, ZN => n3077);
   U2158 : OAI22_X1 port map( A1 => n9309, A2 => n9559, B1 => n8486, B2 => 
                           n9566, ZN => n3078);
   U2159 : OAI22_X1 port map( A1 => n9306, A2 => n9559, B1 => n8487, B2 => 
                           n9566, ZN => n3079);
   U2160 : OAI22_X1 port map( A1 => n9303, A2 => n9559, B1 => n8488, B2 => 
                           n9566, ZN => n3080);
   U2161 : OAI22_X1 port map( A1 => n9300, A2 => n9559, B1 => n8489, B2 => 
                           n9566, ZN => n3081);
   U2162 : OAI22_X1 port map( A1 => n9297, A2 => n9560, B1 => n8490, B2 => 
                           n9565, ZN => n3082);
   U2163 : OAI22_X1 port map( A1 => n9294, A2 => n9560, B1 => n8491, B2 => 
                           n9565, ZN => n3083);
   U2164 : OAI22_X1 port map( A1 => n9291, A2 => n9560, B1 => n8492, B2 => 
                           n9565, ZN => n3084);
   U2165 : OAI22_X1 port map( A1 => n9288, A2 => n9560, B1 => n8493, B2 => 
                           n9565, ZN => n3085);
   U2166 : OAI22_X1 port map( A1 => n9285, A2 => n9560, B1 => n8494, B2 => 
                           n9564, ZN => n3086);
   U2167 : OAI22_X1 port map( A1 => n9282, A2 => n9560, B1 => n8495, B2 => 
                           n9564, ZN => n3087);
   U2168 : OAI22_X1 port map( A1 => n9279, A2 => n9560, B1 => n8496, B2 => 
                           n9564, ZN => n3088);
   U2169 : OAI22_X1 port map( A1 => n9276, A2 => n9560, B1 => n8497, B2 => 
                           n9564, ZN => n3089);
   U2170 : OAI22_X1 port map( A1 => n9273, A2 => n9560, B1 => n8498, B2 => 
                           n9563, ZN => n3090);
   U2171 : OAI22_X1 port map( A1 => n9270, A2 => n9560, B1 => n8499, B2 => 
                           n9563, ZN => n3091);
   U2172 : OAI22_X1 port map( A1 => n9267, A2 => n9560, B1 => n8500, B2 => 
                           n9563, ZN => n3092);
   U2173 : OAI22_X1 port map( A1 => n9264, A2 => n9560, B1 => n8501, B2 => 
                           n9563, ZN => n3093);
   U2174 : OAI22_X1 port map( A1 => n9261, A2 => n9559, B1 => n8502, B2 => 
                           n9562, ZN => n3094);
   U2175 : OAI22_X1 port map( A1 => n9258, A2 => n9560, B1 => n8503, B2 => 
                           n9562, ZN => n3095);
   U2176 : OAI22_X1 port map( A1 => n9255, A2 => n9559, B1 => n8504, B2 => 
                           n9562, ZN => n3096);
   U2177 : OAI22_X1 port map( A1 => n9252, A2 => n9560, B1 => n8505, B2 => 
                           n9562, ZN => n3097);
   U2178 : OAI22_X1 port map( A1 => n9249, A2 => n9559, B1 => n8506, B2 => 
                           n9561, ZN => n3098);
   U2179 : OAI22_X1 port map( A1 => n9246, A2 => n9560, B1 => n8507, B2 => 
                           n9561, ZN => n3099);
   U2180 : OAI22_X1 port map( A1 => n9243, A2 => n9559, B1 => n8508, B2 => 
                           n9561, ZN => n3100);
   U2181 : OAI22_X1 port map( A1 => n9240, A2 => n9560, B1 => n8509, B2 => 
                           n9561, ZN => n3101);
   U2182 : OAI22_X1 port map( A1 => n9330, A2 => n9581, B1 => n8567, B2 => 
                           n9590, ZN => n3135);
   U2183 : OAI22_X1 port map( A1 => n9327, A2 => n9581, B1 => n8568, B2 => 
                           n9590, ZN => n3136);
   U2184 : OAI22_X1 port map( A1 => n9324, A2 => n9581, B1 => n8569, B2 => 
                           n9590, ZN => n3137);
   U2185 : OAI22_X1 port map( A1 => n9321, A2 => n9581, B1 => n8570, B2 => 
                           n9589, ZN => n3138);
   U2186 : OAI22_X1 port map( A1 => n9318, A2 => n9581, B1 => n8571, B2 => 
                           n9589, ZN => n3139);
   U2187 : OAI22_X1 port map( A1 => n9315, A2 => n9581, B1 => n8572, B2 => 
                           n9589, ZN => n3140);
   U2188 : OAI22_X1 port map( A1 => n9312, A2 => n9581, B1 => n8573, B2 => 
                           n9589, ZN => n3141);
   U2189 : OAI22_X1 port map( A1 => n9309, A2 => n9581, B1 => n8574, B2 => 
                           n9588, ZN => n3142);
   U2190 : OAI22_X1 port map( A1 => n9306, A2 => n9581, B1 => n8575, B2 => 
                           n9588, ZN => n3143);
   U2191 : OAI22_X1 port map( A1 => n9303, A2 => n9581, B1 => n8576, B2 => 
                           n9588, ZN => n3144);
   U2192 : OAI22_X1 port map( A1 => n9300, A2 => n9581, B1 => n8577, B2 => 
                           n9588, ZN => n3145);
   U2193 : OAI22_X1 port map( A1 => n9297, A2 => n9582, B1 => n8578, B2 => 
                           n9587, ZN => n3146);
   U2194 : OAI22_X1 port map( A1 => n9294, A2 => n9582, B1 => n8579, B2 => 
                           n9587, ZN => n3147);
   U2195 : OAI22_X1 port map( A1 => n9291, A2 => n9582, B1 => n8580, B2 => 
                           n9587, ZN => n3148);
   U2196 : OAI22_X1 port map( A1 => n9288, A2 => n9582, B1 => n8581, B2 => 
                           n9587, ZN => n3149);
   U2197 : OAI22_X1 port map( A1 => n9285, A2 => n9582, B1 => n8582, B2 => 
                           n9586, ZN => n3150);
   U2198 : OAI22_X1 port map( A1 => n9282, A2 => n9582, B1 => n8583, B2 => 
                           n9586, ZN => n3151);
   U2199 : OAI22_X1 port map( A1 => n9279, A2 => n9582, B1 => n8584, B2 => 
                           n9586, ZN => n3152);
   U2200 : OAI22_X1 port map( A1 => n9276, A2 => n9582, B1 => n8585, B2 => 
                           n9586, ZN => n3153);
   U2201 : OAI22_X1 port map( A1 => n9273, A2 => n9582, B1 => n8586, B2 => 
                           n9585, ZN => n3154);
   U2202 : OAI22_X1 port map( A1 => n9270, A2 => n9582, B1 => n8587, B2 => 
                           n9585, ZN => n3155);
   U2203 : OAI22_X1 port map( A1 => n9267, A2 => n9582, B1 => n8588, B2 => 
                           n9585, ZN => n3156);
   U2204 : OAI22_X1 port map( A1 => n9264, A2 => n9582, B1 => n8589, B2 => 
                           n9585, ZN => n3157);
   U2205 : OAI22_X1 port map( A1 => n9261, A2 => n9581, B1 => n8590, B2 => 
                           n9584, ZN => n3158);
   U2206 : OAI22_X1 port map( A1 => n9258, A2 => n9582, B1 => n8591, B2 => 
                           n9584, ZN => n3159);
   U2207 : OAI22_X1 port map( A1 => n9255, A2 => n9581, B1 => n8592, B2 => 
                           n9584, ZN => n3160);
   U2208 : OAI22_X1 port map( A1 => n9252, A2 => n9582, B1 => n8593, B2 => 
                           n9584, ZN => n3161);
   U2209 : OAI22_X1 port map( A1 => n9249, A2 => n9581, B1 => n8594, B2 => 
                           n9583, ZN => n3162);
   U2210 : OAI22_X1 port map( A1 => n9246, A2 => n9582, B1 => n8595, B2 => 
                           n9583, ZN => n3163);
   U2211 : OAI22_X1 port map( A1 => n9243, A2 => n9581, B1 => n8596, B2 => 
                           n9583, ZN => n3164);
   U2212 : OAI22_X1 port map( A1 => n9240, A2 => n9582, B1 => n8597, B2 => 
                           n9583, ZN => n3165);
   U2213 : OAI22_X1 port map( A1 => n9329, A2 => n9636, B1 => n8775, B2 => 
                           n9645, ZN => n3295);
   U2214 : OAI22_X1 port map( A1 => n9326, A2 => n9636, B1 => n8776, B2 => 
                           n9645, ZN => n3296);
   U2215 : OAI22_X1 port map( A1 => n9323, A2 => n9636, B1 => n8777, B2 => 
                           n9645, ZN => n3297);
   U2216 : OAI22_X1 port map( A1 => n9320, A2 => n9636, B1 => n8778, B2 => 
                           n9644, ZN => n3298);
   U2217 : OAI22_X1 port map( A1 => n9317, A2 => n9636, B1 => n8779, B2 => 
                           n9644, ZN => n3299);
   U2218 : OAI22_X1 port map( A1 => n9311, A2 => n9636, B1 => n8781, B2 => 
                           n9644, ZN => n3301);
   U2219 : OAI22_X1 port map( A1 => n9308, A2 => n9636, B1 => n8782, B2 => 
                           n9643, ZN => n3302);
   U2220 : OAI22_X1 port map( A1 => n9305, A2 => n9636, B1 => n8783, B2 => 
                           n9643, ZN => n3303);
   U2221 : OAI22_X1 port map( A1 => n9302, A2 => n9636, B1 => n8784, B2 => 
                           n9643, ZN => n3304);
   U2222 : OAI22_X1 port map( A1 => n9299, A2 => n9636, B1 => n8785, B2 => 
                           n9643, ZN => n3305);
   U2223 : OAI22_X1 port map( A1 => n9296, A2 => n9637, B1 => n8786, B2 => 
                           n9642, ZN => n3306);
   U2224 : OAI22_X1 port map( A1 => n9290, A2 => n9637, B1 => n8788, B2 => 
                           n9642, ZN => n3308);
   U2225 : OAI22_X1 port map( A1 => n9287, A2 => n9637, B1 => n8789, B2 => 
                           n9642, ZN => n3309);
   U2226 : OAI22_X1 port map( A1 => n9284, A2 => n9637, B1 => n8790, B2 => 
                           n9641, ZN => n3310);
   U2227 : OAI22_X1 port map( A1 => n9278, A2 => n9637, B1 => n8792, B2 => 
                           n9641, ZN => n3312);
   U2228 : OAI22_X1 port map( A1 => n9275, A2 => n9637, B1 => n8793, B2 => 
                           n9641, ZN => n3313);
   U2229 : OAI22_X1 port map( A1 => n9272, A2 => n9637, B1 => n8794, B2 => 
                           n9640, ZN => n3314);
   U2230 : OAI22_X1 port map( A1 => n9269, A2 => n9637, B1 => n8795, B2 => 
                           n9640, ZN => n3315);
   U2231 : OAI22_X1 port map( A1 => n9266, A2 => n9637, B1 => n8796, B2 => 
                           n9640, ZN => n3316);
   U2232 : OAI22_X1 port map( A1 => n9263, A2 => n9637, B1 => n8797, B2 => 
                           n9640, ZN => n3317);
   U2233 : OAI22_X1 port map( A1 => n9332, A2 => n9647, B1 => n8798, B2 => 
                           n9656, ZN => n3326);
   U2234 : OAI22_X1 port map( A1 => n9329, A2 => n9647, B1 => n8799, B2 => 
                           n9656, ZN => n3327);
   U2235 : OAI22_X1 port map( A1 => n9326, A2 => n9647, B1 => n8800, B2 => 
                           n9656, ZN => n3328);
   U2236 : OAI22_X1 port map( A1 => n9323, A2 => n9647, B1 => n8801, B2 => 
                           n9656, ZN => n3329);
   U2237 : OAI22_X1 port map( A1 => n9320, A2 => n9647, B1 => n8802, B2 => 
                           n9655, ZN => n3330);
   U2238 : OAI22_X1 port map( A1 => n9317, A2 => n9647, B1 => n8803, B2 => 
                           n9655, ZN => n3331);
   U2239 : OAI22_X1 port map( A1 => n9314, A2 => n9647, B1 => n8804, B2 => 
                           n9655, ZN => n3332);
   U2240 : OAI22_X1 port map( A1 => n9311, A2 => n9647, B1 => n8805, B2 => 
                           n9655, ZN => n3333);
   U2241 : OAI22_X1 port map( A1 => n9308, A2 => n9647, B1 => n8806, B2 => 
                           n9654, ZN => n3334);
   U2242 : OAI22_X1 port map( A1 => n9305, A2 => n9647, B1 => n8807, B2 => 
                           n9654, ZN => n3335);
   U2243 : OAI22_X1 port map( A1 => n9302, A2 => n9647, B1 => n8808, B2 => 
                           n9654, ZN => n3336);
   U2244 : OAI22_X1 port map( A1 => n9299, A2 => n9647, B1 => n8809, B2 => 
                           n9654, ZN => n3337);
   U2245 : OAI22_X1 port map( A1 => n9296, A2 => n9648, B1 => n8810, B2 => 
                           n9653, ZN => n3338);
   U2246 : OAI22_X1 port map( A1 => n9293, A2 => n9648, B1 => n8811, B2 => 
                           n9653, ZN => n3339);
   U2247 : OAI22_X1 port map( A1 => n9290, A2 => n9648, B1 => n8812, B2 => 
                           n9653, ZN => n3340);
   U2248 : OAI22_X1 port map( A1 => n9287, A2 => n9648, B1 => n8813, B2 => 
                           n9653, ZN => n3341);
   U2249 : OAI22_X1 port map( A1 => n9284, A2 => n9648, B1 => n8814, B2 => 
                           n9652, ZN => n3342);
   U2250 : OAI22_X1 port map( A1 => n9281, A2 => n9648, B1 => n8815, B2 => 
                           n9652, ZN => n3343);
   U2251 : OAI22_X1 port map( A1 => n9278, A2 => n9648, B1 => n8816, B2 => 
                           n9652, ZN => n3344);
   U2252 : OAI22_X1 port map( A1 => n9275, A2 => n9648, B1 => n8817, B2 => 
                           n9652, ZN => n3345);
   U2253 : OAI22_X1 port map( A1 => n9272, A2 => n9648, B1 => n8818, B2 => 
                           n9651, ZN => n3346);
   U2254 : OAI22_X1 port map( A1 => n9269, A2 => n9648, B1 => n8819, B2 => 
                           n9651, ZN => n3347);
   U2255 : OAI22_X1 port map( A1 => n9266, A2 => n9648, B1 => n8820, B2 => 
                           n9651, ZN => n3348);
   U2256 : OAI22_X1 port map( A1 => n9263, A2 => n9648, B1 => n8821, B2 => 
                           n9651, ZN => n3349);
   U2257 : OAI22_X1 port map( A1 => n9260, A2 => n9647, B1 => n8822, B2 => 
                           n9650, ZN => n3350);
   U2258 : OAI22_X1 port map( A1 => n9257, A2 => n9648, B1 => n8823, B2 => 
                           n9650, ZN => n3351);
   U2259 : OAI22_X1 port map( A1 => n9254, A2 => n9647, B1 => n8824, B2 => 
                           n9650, ZN => n3352);
   U2260 : OAI22_X1 port map( A1 => n9251, A2 => n9648, B1 => n8825, B2 => 
                           n9650, ZN => n3353);
   U2261 : OAI22_X1 port map( A1 => n9248, A2 => n9647, B1 => n8826, B2 => 
                           n9649, ZN => n3354);
   U2262 : OAI22_X1 port map( A1 => n9245, A2 => n9648, B1 => n8827, B2 => 
                           n9649, ZN => n3355);
   U2263 : OAI22_X1 port map( A1 => n9242, A2 => n9647, B1 => n8828, B2 => 
                           n9649, ZN => n3356);
   U2264 : OAI22_X1 port map( A1 => n9239, A2 => n9648, B1 => n8829, B2 => 
                           n9649, ZN => n3357);
   U2265 : OAI22_X1 port map( A1 => n9332, A2 => n9669, B1 => n8886, B2 => 
                           n9678, ZN => n3390);
   U2266 : OAI22_X1 port map( A1 => n9329, A2 => n9669, B1 => n8887, B2 => 
                           n9678, ZN => n3391);
   U2267 : OAI22_X1 port map( A1 => n9326, A2 => n9669, B1 => n8888, B2 => 
                           n9678, ZN => n3392);
   U2268 : OAI22_X1 port map( A1 => n9323, A2 => n9669, B1 => n8889, B2 => 
                           n9678, ZN => n3393);
   U2269 : OAI22_X1 port map( A1 => n9320, A2 => n9669, B1 => n8890, B2 => 
                           n9677, ZN => n3394);
   U2270 : OAI22_X1 port map( A1 => n9317, A2 => n9669, B1 => n8891, B2 => 
                           n9677, ZN => n3395);
   U2271 : OAI22_X1 port map( A1 => n9314, A2 => n9669, B1 => n8892, B2 => 
                           n9677, ZN => n3396);
   U2272 : OAI22_X1 port map( A1 => n9311, A2 => n9669, B1 => n8893, B2 => 
                           n9677, ZN => n3397);
   U2273 : OAI22_X1 port map( A1 => n9308, A2 => n9669, B1 => n8894, B2 => 
                           n9676, ZN => n3398);
   U2274 : OAI22_X1 port map( A1 => n9305, A2 => n9669, B1 => n8895, B2 => 
                           n9676, ZN => n3399);
   U2275 : OAI22_X1 port map( A1 => n9302, A2 => n9669, B1 => n8896, B2 => 
                           n9676, ZN => n3400);
   U2276 : OAI22_X1 port map( A1 => n9299, A2 => n9669, B1 => n8897, B2 => 
                           n9676, ZN => n3401);
   U2277 : OAI22_X1 port map( A1 => n9296, A2 => n9670, B1 => n8898, B2 => 
                           n9675, ZN => n3402);
   U2278 : OAI22_X1 port map( A1 => n9293, A2 => n9670, B1 => n8899, B2 => 
                           n9675, ZN => n3403);
   U2279 : OAI22_X1 port map( A1 => n9290, A2 => n9670, B1 => n8900, B2 => 
                           n9675, ZN => n3404);
   U2280 : OAI22_X1 port map( A1 => n9287, A2 => n9670, B1 => n8901, B2 => 
                           n9675, ZN => n3405);
   U2281 : OAI22_X1 port map( A1 => n9284, A2 => n9670, B1 => n8902, B2 => 
                           n9674, ZN => n3406);
   U2282 : OAI22_X1 port map( A1 => n9281, A2 => n9670, B1 => n8903, B2 => 
                           n9674, ZN => n3407);
   U2283 : OAI22_X1 port map( A1 => n9278, A2 => n9670, B1 => n8904, B2 => 
                           n9674, ZN => n3408);
   U2284 : OAI22_X1 port map( A1 => n9275, A2 => n9670, B1 => n8905, B2 => 
                           n9674, ZN => n3409);
   U2285 : OAI22_X1 port map( A1 => n9272, A2 => n9670, B1 => n8906, B2 => 
                           n9673, ZN => n3410);
   U2286 : OAI22_X1 port map( A1 => n9269, A2 => n9670, B1 => n8907, B2 => 
                           n9673, ZN => n3411);
   U2287 : OAI22_X1 port map( A1 => n9266, A2 => n9670, B1 => n8908, B2 => 
                           n9673, ZN => n3412);
   U2288 : OAI22_X1 port map( A1 => n9263, A2 => n9670, B1 => n8909, B2 => 
                           n9673, ZN => n3413);
   U2289 : OAI22_X1 port map( A1 => n9260, A2 => n9669, B1 => n8910, B2 => 
                           n9672, ZN => n3414);
   U2290 : OAI22_X1 port map( A1 => n9257, A2 => n9670, B1 => n8911, B2 => 
                           n9672, ZN => n3415);
   U2291 : OAI22_X1 port map( A1 => n9254, A2 => n9669, B1 => n8912, B2 => 
                           n9672, ZN => n3416);
   U2292 : OAI22_X1 port map( A1 => n9251, A2 => n9670, B1 => n8913, B2 => 
                           n9672, ZN => n3417);
   U2293 : OAI22_X1 port map( A1 => n9248, A2 => n9669, B1 => n8914, B2 => 
                           n9671, ZN => n3418);
   U2294 : OAI22_X1 port map( A1 => n9245, A2 => n9670, B1 => n8915, B2 => 
                           n9671, ZN => n3419);
   U2295 : OAI22_X1 port map( A1 => n9242, A2 => n9669, B1 => n8916, B2 => 
                           n9671, ZN => n3420);
   U2296 : OAI22_X1 port map( A1 => n9239, A2 => n9670, B1 => n8917, B2 => 
                           n9671, ZN => n3421);
   U2297 : OAI22_X1 port map( A1 => n9331, A2 => n9846, B1 => n8244, B2 => 
                           n9847, ZN => n9141);
   U2298 : OAI22_X1 port map( A1 => n9328, A2 => n9845, B1 => n8242, B2 => 
                           n9847, ZN => n9140);
   U2299 : OAI22_X1 port map( A1 => n9325, A2 => n9846, B1 => n8240, B2 => 
                           n9847, ZN => n9139);
   U2300 : OAI22_X1 port map( A1 => n9322, A2 => n9845, B1 => n8238, B2 => 
                           n9847, ZN => n9138);
   U2301 : OAI22_X1 port map( A1 => n9319, A2 => n9846, B1 => n8236, B2 => 
                           n9848, ZN => n9137);
   U2302 : OAI22_X1 port map( A1 => n9316, A2 => n9845, B1 => n8234, B2 => 
                           n9848, ZN => n9136);
   U2303 : OAI22_X1 port map( A1 => n9313, A2 => n9846, B1 => n8232, B2 => 
                           n9848, ZN => n9135);
   U2304 : OAI22_X1 port map( A1 => n9310, A2 => n9845, B1 => n8230, B2 => 
                           n9848, ZN => n9134);
   U2305 : OAI22_X1 port map( A1 => n9307, A2 => n9846, B1 => n8228, B2 => 
                           n9849, ZN => n9133);
   U2306 : OAI22_X1 port map( A1 => n9304, A2 => n9846, B1 => n8226, B2 => 
                           n9849, ZN => n9132);
   U2307 : OAI22_X1 port map( A1 => n9301, A2 => n9846, B1 => n8224, B2 => 
                           n9849, ZN => n9131);
   U2308 : OAI22_X1 port map( A1 => n9298, A2 => n9846, B1 => n8222, B2 => 
                           n9849, ZN => n9130);
   U2309 : OAI22_X1 port map( A1 => n9295, A2 => n9846, B1 => n8220, B2 => 
                           n9850, ZN => n9129);
   U2310 : OAI22_X1 port map( A1 => n9292, A2 => n9846, B1 => n8218, B2 => 
                           n9850, ZN => n9128);
   U2311 : OAI22_X1 port map( A1 => n9289, A2 => n9846, B1 => n8216, B2 => 
                           n9850, ZN => n9127);
   U2312 : OAI22_X1 port map( A1 => n9286, A2 => n9846, B1 => n8214, B2 => 
                           n9850, ZN => n9126);
   U2313 : OAI22_X1 port map( A1 => n9283, A2 => n9846, B1 => n8212, B2 => 
                           n9851, ZN => n9125);
   U2314 : OAI22_X1 port map( A1 => n9280, A2 => n9846, B1 => n8210, B2 => 
                           n9851, ZN => n9124);
   U2315 : OAI22_X1 port map( A1 => n9277, A2 => n9846, B1 => n8208, B2 => 
                           n9851, ZN => n9123);
   U2316 : OAI22_X1 port map( A1 => n9274, A2 => n9846, B1 => n8206, B2 => 
                           n9851, ZN => n9122);
   U2317 : OAI22_X1 port map( A1 => n9271, A2 => n9845, B1 => n8204, B2 => 
                           n9852, ZN => n9121);
   U2318 : OAI22_X1 port map( A1 => n9268, A2 => n9845, B1 => n8202, B2 => 
                           n9852, ZN => n9120);
   U2319 : OAI22_X1 port map( A1 => n9265, A2 => n9845, B1 => n8200, B2 => 
                           n9852, ZN => n9119);
   U2320 : OAI22_X1 port map( A1 => n9262, A2 => n9845, B1 => n8198, B2 => 
                           n9852, ZN => n9118);
   U2321 : OAI22_X1 port map( A1 => n9260, A2 => n9614, B1 => n8287, B2 => 
                           n9617, ZN => n3254);
   U2322 : OAI22_X1 port map( A1 => n9257, A2 => n9615, B1 => n8288, B2 => 
                           n9617, ZN => n3255);
   U2323 : OAI22_X1 port map( A1 => n9254, A2 => n9614, B1 => n8289, B2 => 
                           n9617, ZN => n3256);
   U2324 : OAI22_X1 port map( A1 => n9251, A2 => n9615, B1 => n8290, B2 => 
                           n9617, ZN => n3257);
   U2325 : OAI22_X1 port map( A1 => n9248, A2 => n9614, B1 => n8291, B2 => 
                           n9616, ZN => n3258);
   U2326 : OAI22_X1 port map( A1 => n9245, A2 => n9615, B1 => n8292, B2 => 
                           n9616, ZN => n3259);
   U2327 : OAI22_X1 port map( A1 => n9242, A2 => n9614, B1 => n8293, B2 => 
                           n9616, ZN => n3260);
   U2328 : OAI22_X1 port map( A1 => n9239, A2 => n9615, B1 => n8294, B2 => 
                           n9616, ZN => n3261);
   U2329 : OAI22_X1 port map( A1 => n9260, A2 => n9658, B1 => n8303, B2 => 
                           n9661, ZN => n3382);
   U2330 : OAI22_X1 port map( A1 => n9257, A2 => n9659, B1 => n8304, B2 => 
                           n9661, ZN => n3383);
   U2331 : OAI22_X1 port map( A1 => n9254, A2 => n9658, B1 => n8305, B2 => 
                           n9661, ZN => n3384);
   U2332 : OAI22_X1 port map( A1 => n9251, A2 => n9659, B1 => n8306, B2 => 
                           n9661, ZN => n3385);
   U2333 : OAI22_X1 port map( A1 => n9248, A2 => n9658, B1 => n8307, B2 => 
                           n9660, ZN => n3386);
   U2334 : OAI22_X1 port map( A1 => n9245, A2 => n9659, B1 => n8308, B2 => 
                           n9660, ZN => n3387);
   U2335 : OAI22_X1 port map( A1 => n9242, A2 => n9658, B1 => n8309, B2 => 
                           n9660, ZN => n3388);
   U2336 : OAI22_X1 port map( A1 => n9239, A2 => n9659, B1 => n8310, B2 => 
                           n9660, ZN => n3389);
   U2337 : OAI22_X1 port map( A1 => n9261, A2 => n9570, B1 => n8319, B2 => 
                           n9573, ZN => n3126);
   U2338 : OAI22_X1 port map( A1 => n9258, A2 => n9571, B1 => n8320, B2 => 
                           n9573, ZN => n3127);
   U2339 : OAI22_X1 port map( A1 => n9255, A2 => n9570, B1 => n8321, B2 => 
                           n9573, ZN => n3128);
   U2340 : OAI22_X1 port map( A1 => n9252, A2 => n9571, B1 => n8322, B2 => 
                           n9573, ZN => n3129);
   U2341 : OAI22_X1 port map( A1 => n9249, A2 => n9570, B1 => n8323, B2 => 
                           n9572, ZN => n3130);
   U2342 : OAI22_X1 port map( A1 => n9246, A2 => n9571, B1 => n8324, B2 => 
                           n9572, ZN => n3131);
   U2343 : OAI22_X1 port map( A1 => n9243, A2 => n9570, B1 => n8325, B2 => 
                           n9572, ZN => n3132);
   U2344 : OAI22_X1 port map( A1 => n9240, A2 => n9571, B1 => n8326, B2 => 
                           n9572, ZN => n3133);
   U2345 : OAI22_X1 port map( A1 => n9259, A2 => n9845, B1 => n8196, B2 => 
                           n9853, ZN => n9117);
   U2346 : OAI22_X1 port map( A1 => n9256, A2 => n9845, B1 => n8194, B2 => 
                           n9853, ZN => n9116);
   U2347 : OAI22_X1 port map( A1 => n9253, A2 => n9845, B1 => n8192, B2 => 
                           n9853, ZN => n9115);
   U2348 : OAI22_X1 port map( A1 => n9250, A2 => n9845, B1 => n8190, B2 => 
                           n9853, ZN => n9114);
   U2349 : OAI22_X1 port map( A1 => n9247, A2 => n9845, B1 => n8188, B2 => 
                           n9854, ZN => n9113);
   U2350 : OAI22_X1 port map( A1 => n9244, A2 => n9845, B1 => n8186, B2 => 
                           n9854, ZN => n9112);
   U2351 : OAI22_X1 port map( A1 => n9241, A2 => n9845, B1 => n8184, B2 => 
                           n9854, ZN => n9111);
   U2352 : OAI22_X1 port map( A1 => n9238, A2 => n9845, B1 => n8182, B2 => 
                           n9854, ZN => n9110);
   U2353 : OAI22_X1 port map( A1 => n9331, A2 => n9780, B1 => n8343, B2 => 
                           n9781, ZN => n3958);
   U2354 : OAI22_X1 port map( A1 => n9328, A2 => n9779, B1 => n8344, B2 => 
                           n9781, ZN => n3942);
   U2355 : OAI22_X1 port map( A1 => n9325, A2 => n9780, B1 => n8345, B2 => 
                           n9781, ZN => n3926);
   U2356 : OAI22_X1 port map( A1 => n9322, A2 => n9779, B1 => n8346, B2 => 
                           n9781, ZN => n3910);
   U2357 : OAI22_X1 port map( A1 => n9319, A2 => n9780, B1 => n8347, B2 => 
                           n9782, ZN => n3894);
   U2358 : OAI22_X1 port map( A1 => n9316, A2 => n9779, B1 => n8348, B2 => 
                           n9782, ZN => n3878);
   U2359 : OAI22_X1 port map( A1 => n9313, A2 => n9780, B1 => n8349, B2 => 
                           n9782, ZN => n3862);
   U2360 : OAI22_X1 port map( A1 => n9310, A2 => n9779, B1 => n8350, B2 => 
                           n9782, ZN => n3846);
   U2361 : OAI22_X1 port map( A1 => n9307, A2 => n9780, B1 => n8351, B2 => 
                           n9783, ZN => n3830);
   U2362 : OAI22_X1 port map( A1 => n9304, A2 => n9780, B1 => n8352, B2 => 
                           n9783, ZN => n3814);
   U2363 : OAI22_X1 port map( A1 => n9301, A2 => n9780, B1 => n8353, B2 => 
                           n9783, ZN => n3798);
   U2364 : OAI22_X1 port map( A1 => n9298, A2 => n9780, B1 => n8354, B2 => 
                           n9783, ZN => n3782);
   U2365 : OAI22_X1 port map( A1 => n9295, A2 => n9780, B1 => n8355, B2 => 
                           n9784, ZN => n3766);
   U2366 : OAI22_X1 port map( A1 => n9292, A2 => n9780, B1 => n8356, B2 => 
                           n9784, ZN => n3750);
   U2367 : OAI22_X1 port map( A1 => n9289, A2 => n9780, B1 => n8357, B2 => 
                           n9784, ZN => n3734);
   U2368 : OAI22_X1 port map( A1 => n9286, A2 => n9780, B1 => n8358, B2 => 
                           n9784, ZN => n3718);
   U2369 : OAI22_X1 port map( A1 => n9283, A2 => n9780, B1 => n8359, B2 => 
                           n9785, ZN => n3702);
   U2370 : OAI22_X1 port map( A1 => n9280, A2 => n9780, B1 => n8360, B2 => 
                           n9785, ZN => n3686);
   U2371 : OAI22_X1 port map( A1 => n9277, A2 => n9780, B1 => n8361, B2 => 
                           n9785, ZN => n3670);
   U2372 : OAI22_X1 port map( A1 => n9274, A2 => n9780, B1 => n8362, B2 => 
                           n9785, ZN => n3654);
   U2373 : OAI22_X1 port map( A1 => n9271, A2 => n9779, B1 => n8363, B2 => 
                           n9786, ZN => n3638);
   U2374 : OAI22_X1 port map( A1 => n9268, A2 => n9779, B1 => n8364, B2 => 
                           n9786, ZN => n3622);
   U2375 : OAI22_X1 port map( A1 => n9265, A2 => n9779, B1 => n8365, B2 => 
                           n9786, ZN => n3606);
   U2376 : OAI22_X1 port map( A1 => n9262, A2 => n9779, B1 => n8366, B2 => 
                           n9786, ZN => n3590);
   U2377 : OAI22_X1 port map( A1 => n9259, A2 => n9779, B1 => n8367, B2 => 
                           n9787, ZN => n3574);
   U2378 : OAI22_X1 port map( A1 => n9256, A2 => n9779, B1 => n8368, B2 => 
                           n9787, ZN => n3558);
   U2379 : OAI22_X1 port map( A1 => n9253, A2 => n9779, B1 => n8369, B2 => 
                           n9787, ZN => n3542);
   U2380 : OAI22_X1 port map( A1 => n9250, A2 => n9779, B1 => n8370, B2 => 
                           n9787, ZN => n3526);
   U2381 : OAI22_X1 port map( A1 => n9247, A2 => n9779, B1 => n8371, B2 => 
                           n9788, ZN => n3510);
   U2382 : OAI22_X1 port map( A1 => n9244, A2 => n9779, B1 => n8372, B2 => 
                           n9788, ZN => n3494);
   U2383 : OAI22_X1 port map( A1 => n9241, A2 => n9779, B1 => n8373, B2 => 
                           n9788, ZN => n3478);
   U2384 : OAI22_X1 port map( A1 => n9238, A2 => n9779, B1 => n8374, B2 => 
                           n9788, ZN => n3462);
   U2385 : OAI22_X1 port map( A1 => n9331, A2 => n9758, B1 => n8407, B2 => 
                           n9759, ZN => n3956);
   U2386 : OAI22_X1 port map( A1 => n9328, A2 => n9757, B1 => n8408, B2 => 
                           n9759, ZN => n3940);
   U2387 : OAI22_X1 port map( A1 => n9325, A2 => n9758, B1 => n8409, B2 => 
                           n9759, ZN => n3924);
   U2388 : OAI22_X1 port map( A1 => n9322, A2 => n9757, B1 => n8410, B2 => 
                           n9759, ZN => n3908);
   U2389 : OAI22_X1 port map( A1 => n9319, A2 => n9758, B1 => n8411, B2 => 
                           n9760, ZN => n3892);
   U2390 : OAI22_X1 port map( A1 => n9316, A2 => n9757, B1 => n8412, B2 => 
                           n9760, ZN => n3876);
   U2391 : OAI22_X1 port map( A1 => n9313, A2 => n9758, B1 => n8413, B2 => 
                           n9760, ZN => n3860);
   U2392 : OAI22_X1 port map( A1 => n9310, A2 => n9757, B1 => n8414, B2 => 
                           n9760, ZN => n3844);
   U2393 : OAI22_X1 port map( A1 => n9307, A2 => n9758, B1 => n8415, B2 => 
                           n9761, ZN => n3828);
   U2394 : OAI22_X1 port map( A1 => n9304, A2 => n9758, B1 => n8416, B2 => 
                           n9761, ZN => n3812);
   U2395 : OAI22_X1 port map( A1 => n9301, A2 => n9758, B1 => n8417, B2 => 
                           n9761, ZN => n3796);
   U2396 : OAI22_X1 port map( A1 => n9298, A2 => n9758, B1 => n8418, B2 => 
                           n9761, ZN => n3780);
   U2397 : OAI22_X1 port map( A1 => n9295, A2 => n9758, B1 => n8419, B2 => 
                           n9762, ZN => n3764);
   U2398 : OAI22_X1 port map( A1 => n9292, A2 => n9758, B1 => n8420, B2 => 
                           n9762, ZN => n3748);
   U2399 : OAI22_X1 port map( A1 => n9289, A2 => n9758, B1 => n8421, B2 => 
                           n9762, ZN => n3732);
   U2400 : OAI22_X1 port map( A1 => n9286, A2 => n9758, B1 => n8422, B2 => 
                           n9762, ZN => n3716);
   U2401 : OAI22_X1 port map( A1 => n9283, A2 => n9758, B1 => n8423, B2 => 
                           n9763, ZN => n3700);
   U2402 : OAI22_X1 port map( A1 => n9280, A2 => n9758, B1 => n8424, B2 => 
                           n9763, ZN => n3684);
   U2403 : OAI22_X1 port map( A1 => n9277, A2 => n9758, B1 => n8425, B2 => 
                           n9763, ZN => n3668);
   U2404 : OAI22_X1 port map( A1 => n9274, A2 => n9758, B1 => n8426, B2 => 
                           n9763, ZN => n3652);
   U2405 : OAI22_X1 port map( A1 => n9271, A2 => n9757, B1 => n8427, B2 => 
                           n9764, ZN => n3636);
   U2406 : OAI22_X1 port map( A1 => n9268, A2 => n9757, B1 => n8428, B2 => 
                           n9764, ZN => n3620);
   U2407 : OAI22_X1 port map( A1 => n9265, A2 => n9757, B1 => n8429, B2 => 
                           n9764, ZN => n3604);
   U2408 : OAI22_X1 port map( A1 => n9262, A2 => n9757, B1 => n8430, B2 => 
                           n9764, ZN => n3588);
   U2409 : OAI22_X1 port map( A1 => n9259, A2 => n9757, B1 => n8431, B2 => 
                           n9765, ZN => n3572);
   U2410 : OAI22_X1 port map( A1 => n9256, A2 => n9757, B1 => n8432, B2 => 
                           n9765, ZN => n3556);
   U2411 : OAI22_X1 port map( A1 => n9253, A2 => n9757, B1 => n8433, B2 => 
                           n9765, ZN => n3540);
   U2412 : OAI22_X1 port map( A1 => n9250, A2 => n9757, B1 => n8434, B2 => 
                           n9765, ZN => n3524);
   U2413 : OAI22_X1 port map( A1 => n9247, A2 => n9757, B1 => n8435, B2 => 
                           n9766, ZN => n3508);
   U2414 : OAI22_X1 port map( A1 => n9244, A2 => n9757, B1 => n8436, B2 => 
                           n9766, ZN => n3492);
   U2415 : OAI22_X1 port map( A1 => n9241, A2 => n9757, B1 => n8437, B2 => 
                           n9766, ZN => n3476);
   U2416 : OAI22_X1 port map( A1 => n9238, A2 => n9757, B1 => n8438, B2 => 
                           n9766, ZN => n3460);
   U2417 : OAI22_X1 port map( A1 => n9333, A2 => n9570, B1 => n8542, B2 => 
                           n9579, ZN => n3102);
   U2418 : OAI22_X1 port map( A1 => n9330, A2 => n9570, B1 => n8543, B2 => 
                           n9579, ZN => n3103);
   U2419 : OAI22_X1 port map( A1 => n9327, A2 => n9570, B1 => n8544, B2 => 
                           n9579, ZN => n3104);
   U2420 : OAI22_X1 port map( A1 => n9324, A2 => n9570, B1 => n8545, B2 => 
                           n9579, ZN => n3105);
   U2421 : OAI22_X1 port map( A1 => n9321, A2 => n9570, B1 => n8546, B2 => 
                           n9578, ZN => n3106);
   U2422 : OAI22_X1 port map( A1 => n9318, A2 => n9570, B1 => n8547, B2 => 
                           n9578, ZN => n3107);
   U2423 : OAI22_X1 port map( A1 => n9315, A2 => n9570, B1 => n8548, B2 => 
                           n9578, ZN => n3108);
   U2424 : OAI22_X1 port map( A1 => n9312, A2 => n9570, B1 => n8549, B2 => 
                           n9578, ZN => n3109);
   U2425 : OAI22_X1 port map( A1 => n9309, A2 => n9570, B1 => n8550, B2 => 
                           n9577, ZN => n3110);
   U2426 : OAI22_X1 port map( A1 => n9306, A2 => n9570, B1 => n8551, B2 => 
                           n9577, ZN => n3111);
   U2427 : OAI22_X1 port map( A1 => n9303, A2 => n9570, B1 => n8552, B2 => 
                           n9577, ZN => n3112);
   U2428 : OAI22_X1 port map( A1 => n9300, A2 => n9570, B1 => n8553, B2 => 
                           n9577, ZN => n3113);
   U2429 : OAI22_X1 port map( A1 => n9297, A2 => n9571, B1 => n8554, B2 => 
                           n9576, ZN => n3114);
   U2430 : OAI22_X1 port map( A1 => n9294, A2 => n9571, B1 => n8555, B2 => 
                           n9576, ZN => n3115);
   U2431 : OAI22_X1 port map( A1 => n9291, A2 => n9571, B1 => n8556, B2 => 
                           n9576, ZN => n3116);
   U2432 : OAI22_X1 port map( A1 => n9288, A2 => n9571, B1 => n8557, B2 => 
                           n9576, ZN => n3117);
   U2433 : OAI22_X1 port map( A1 => n9285, A2 => n9571, B1 => n8558, B2 => 
                           n9575, ZN => n3118);
   U2434 : OAI22_X1 port map( A1 => n9282, A2 => n9571, B1 => n8559, B2 => 
                           n9575, ZN => n3119);
   U2435 : OAI22_X1 port map( A1 => n9279, A2 => n9571, B1 => n8560, B2 => 
                           n9575, ZN => n3120);
   U2436 : OAI22_X1 port map( A1 => n9276, A2 => n9571, B1 => n8561, B2 => 
                           n9575, ZN => n3121);
   U2437 : OAI22_X1 port map( A1 => n9273, A2 => n9571, B1 => n8562, B2 => 
                           n9574, ZN => n3122);
   U2438 : OAI22_X1 port map( A1 => n9270, A2 => n9571, B1 => n8563, B2 => 
                           n9574, ZN => n3123);
   U2439 : OAI22_X1 port map( A1 => n9267, A2 => n9571, B1 => n8564, B2 => 
                           n9574, ZN => n3124);
   U2440 : OAI22_X1 port map( A1 => n9264, A2 => n9571, B1 => n8565, B2 => 
                           n9574, ZN => n3125);
   U2441 : OAI22_X1 port map( A1 => n9332, A2 => n9614, B1 => n8718, B2 => 
                           n9623, ZN => n3230);
   U2442 : OAI22_X1 port map( A1 => n9329, A2 => n9614, B1 => n8719, B2 => 
                           n9623, ZN => n3231);
   U2443 : OAI22_X1 port map( A1 => n9326, A2 => n9614, B1 => n8720, B2 => 
                           n9623, ZN => n3232);
   U2444 : OAI22_X1 port map( A1 => n9323, A2 => n9614, B1 => n8721, B2 => 
                           n9623, ZN => n3233);
   U2445 : OAI22_X1 port map( A1 => n9320, A2 => n9614, B1 => n8722, B2 => 
                           n9622, ZN => n3234);
   U2446 : OAI22_X1 port map( A1 => n9317, A2 => n9614, B1 => n8723, B2 => 
                           n9622, ZN => n3235);
   U2447 : OAI22_X1 port map( A1 => n9314, A2 => n9614, B1 => n8724, B2 => 
                           n9622, ZN => n3236);
   U2448 : OAI22_X1 port map( A1 => n9311, A2 => n9614, B1 => n8725, B2 => 
                           n9622, ZN => n3237);
   U2449 : OAI22_X1 port map( A1 => n9308, A2 => n9614, B1 => n8726, B2 => 
                           n9621, ZN => n3238);
   U2450 : OAI22_X1 port map( A1 => n9305, A2 => n9614, B1 => n8727, B2 => 
                           n9621, ZN => n3239);
   U2451 : OAI22_X1 port map( A1 => n9302, A2 => n9614, B1 => n8728, B2 => 
                           n9621, ZN => n3240);
   U2452 : OAI22_X1 port map( A1 => n9299, A2 => n9614, B1 => n8729, B2 => 
                           n9621, ZN => n3241);
   U2453 : OAI22_X1 port map( A1 => n9296, A2 => n9615, B1 => n8730, B2 => 
                           n9620, ZN => n3242);
   U2454 : OAI22_X1 port map( A1 => n9293, A2 => n9615, B1 => n8731, B2 => 
                           n9620, ZN => n3243);
   U2455 : OAI22_X1 port map( A1 => n9290, A2 => n9615, B1 => n8732, B2 => 
                           n9620, ZN => n3244);
   U2456 : OAI22_X1 port map( A1 => n9287, A2 => n9615, B1 => n8733, B2 => 
                           n9620, ZN => n3245);
   U2457 : OAI22_X1 port map( A1 => n9284, A2 => n9615, B1 => n8734, B2 => 
                           n9619, ZN => n3246);
   U2458 : OAI22_X1 port map( A1 => n9281, A2 => n9615, B1 => n8735, B2 => 
                           n9619, ZN => n3247);
   U2459 : OAI22_X1 port map( A1 => n9278, A2 => n9615, B1 => n8736, B2 => 
                           n9619, ZN => n3248);
   U2460 : OAI22_X1 port map( A1 => n9275, A2 => n9615, B1 => n8737, B2 => 
                           n9619, ZN => n3249);
   U2461 : OAI22_X1 port map( A1 => n9272, A2 => n9615, B1 => n8738, B2 => 
                           n9618, ZN => n3250);
   U2462 : OAI22_X1 port map( A1 => n9269, A2 => n9615, B1 => n8739, B2 => 
                           n9618, ZN => n3251);
   U2463 : OAI22_X1 port map( A1 => n9266, A2 => n9615, B1 => n8740, B2 => 
                           n9618, ZN => n3252);
   U2464 : OAI22_X1 port map( A1 => n9263, A2 => n9615, B1 => n8741, B2 => 
                           n9618, ZN => n3253);
   U2465 : OAI22_X1 port map( A1 => n9328, A2 => n9812, B1 => n8243, B2 => 
                           n9821, ZN => n9015);
   U2466 : OAI22_X1 port map( A1 => n9325, A2 => n9812, B1 => n8241, B2 => 
                           n9821, ZN => n9016);
   U2467 : OAI22_X1 port map( A1 => n9322, A2 => n9812, B1 => n8239, B2 => 
                           n9821, ZN => n9017);
   U2468 : OAI22_X1 port map( A1 => n9319, A2 => n9812, B1 => n8237, B2 => 
                           n9820, ZN => n9018);
   U2469 : OAI22_X1 port map( A1 => n9316, A2 => n9812, B1 => n8235, B2 => 
                           n9820, ZN => n9019);
   U2470 : OAI22_X1 port map( A1 => n9310, A2 => n9812, B1 => n8231, B2 => 
                           n9820, ZN => n9021);
   U2471 : OAI22_X1 port map( A1 => n9307, A2 => n9812, B1 => n8229, B2 => 
                           n9819, ZN => n9022);
   U2472 : OAI22_X1 port map( A1 => n9304, A2 => n9812, B1 => n8227, B2 => 
                           n9819, ZN => n9023);
   U2473 : OAI22_X1 port map( A1 => n9301, A2 => n9812, B1 => n8225, B2 => 
                           n9819, ZN => n9024);
   U2474 : OAI22_X1 port map( A1 => n9298, A2 => n9812, B1 => n8223, B2 => 
                           n9819, ZN => n9025);
   U2475 : OAI22_X1 port map( A1 => n9295, A2 => n9813, B1 => n8221, B2 => 
                           n9818, ZN => n9026);
   U2476 : OAI22_X1 port map( A1 => n9289, A2 => n9813, B1 => n8217, B2 => 
                           n9818, ZN => n9028);
   U2477 : OAI22_X1 port map( A1 => n9286, A2 => n9813, B1 => n8215, B2 => 
                           n9818, ZN => n9029);
   U2478 : OAI22_X1 port map( A1 => n9283, A2 => n9813, B1 => n8213, B2 => 
                           n9817, ZN => n9030);
   U2479 : OAI22_X1 port map( A1 => n9277, A2 => n9813, B1 => n8209, B2 => 
                           n9817, ZN => n9032);
   U2480 : OAI22_X1 port map( A1 => n9274, A2 => n9813, B1 => n8207, B2 => 
                           n9817, ZN => n9033);
   U2481 : OAI22_X1 port map( A1 => n9271, A2 => n9813, B1 => n8205, B2 => 
                           n9816, ZN => n9034);
   U2482 : OAI22_X1 port map( A1 => n9268, A2 => n9813, B1 => n8203, B2 => 
                           n9816, ZN => n9035);
   U2483 : OAI22_X1 port map( A1 => n9265, A2 => n9813, B1 => n8201, B2 => 
                           n9816, ZN => n9036);
   U2484 : OAI22_X1 port map( A1 => n9262, A2 => n9813, B1 => n8199, B2 => 
                           n9816, ZN => n9037);
   U2485 : OAI22_X1 port map( A1 => n9259, A2 => n9812, B1 => n8197, B2 => 
                           n9815, ZN => n9038);
   U2486 : OAI22_X1 port map( A1 => n9256, A2 => n9813, B1 => n8195, B2 => 
                           n9815, ZN => n9039);
   U2487 : OAI22_X1 port map( A1 => n9253, A2 => n9812, B1 => n8193, B2 => 
                           n9815, ZN => n9040);
   U2488 : OAI22_X1 port map( A1 => n9250, A2 => n9813, B1 => n8191, B2 => 
                           n9815, ZN => n9041);
   U2489 : OAI22_X1 port map( A1 => n9247, A2 => n9812, B1 => n8189, B2 => 
                           n9814, ZN => n9042);
   U2490 : OAI22_X1 port map( A1 => n9244, A2 => n9813, B1 => n8187, B2 => 
                           n9814, ZN => n9043);
   U2491 : OAI22_X1 port map( A1 => n9241, A2 => n9812, B1 => n8185, B2 => 
                           n9814, ZN => n9044);
   U2492 : OAI22_X1 port map( A1 => n9238, A2 => n9813, B1 => n8183, B2 => 
                           n9814, ZN => n9045);
   U2493 : OAI22_X1 port map( A1 => n9332, A2 => n9658, B1 => n8862, B2 => 
                           n9667, ZN => n3358);
   U2494 : OAI22_X1 port map( A1 => n9329, A2 => n9658, B1 => n8863, B2 => 
                           n9667, ZN => n3359);
   U2495 : OAI22_X1 port map( A1 => n9326, A2 => n9658, B1 => n8864, B2 => 
                           n9667, ZN => n3360);
   U2496 : OAI22_X1 port map( A1 => n9323, A2 => n9658, B1 => n8865, B2 => 
                           n9667, ZN => n3361);
   U2497 : OAI22_X1 port map( A1 => n9320, A2 => n9658, B1 => n8866, B2 => 
                           n9666, ZN => n3362);
   U2498 : OAI22_X1 port map( A1 => n9317, A2 => n9658, B1 => n8867, B2 => 
                           n9666, ZN => n3363);
   U2499 : OAI22_X1 port map( A1 => n9314, A2 => n9658, B1 => n8868, B2 => 
                           n9666, ZN => n3364);
   U2500 : OAI22_X1 port map( A1 => n9311, A2 => n9658, B1 => n8869, B2 => 
                           n9666, ZN => n3365);
   U2501 : OAI22_X1 port map( A1 => n9308, A2 => n9658, B1 => n8870, B2 => 
                           n9665, ZN => n3366);
   U2502 : OAI22_X1 port map( A1 => n9305, A2 => n9658, B1 => n8871, B2 => 
                           n9665, ZN => n3367);
   U2503 : OAI22_X1 port map( A1 => n9302, A2 => n9658, B1 => n8872, B2 => 
                           n9665, ZN => n3368);
   U2504 : OAI22_X1 port map( A1 => n9299, A2 => n9658, B1 => n8873, B2 => 
                           n9665, ZN => n3369);
   U2505 : OAI22_X1 port map( A1 => n9296, A2 => n9659, B1 => n8874, B2 => 
                           n9664, ZN => n3370);
   U2506 : OAI22_X1 port map( A1 => n9293, A2 => n9659, B1 => n8875, B2 => 
                           n9664, ZN => n3371);
   U2507 : OAI22_X1 port map( A1 => n9290, A2 => n9659, B1 => n8876, B2 => 
                           n9664, ZN => n3372);
   U2508 : OAI22_X1 port map( A1 => n9287, A2 => n9659, B1 => n8877, B2 => 
                           n9664, ZN => n3373);
   U2509 : OAI22_X1 port map( A1 => n9284, A2 => n9659, B1 => n8878, B2 => 
                           n9663, ZN => n3374);
   U2510 : OAI22_X1 port map( A1 => n9281, A2 => n9659, B1 => n8879, B2 => 
                           n9663, ZN => n3375);
   U2511 : OAI22_X1 port map( A1 => n9278, A2 => n9659, B1 => n8880, B2 => 
                           n9663, ZN => n3376);
   U2512 : OAI22_X1 port map( A1 => n9275, A2 => n9659, B1 => n8881, B2 => 
                           n9663, ZN => n3377);
   U2513 : OAI22_X1 port map( A1 => n9272, A2 => n9659, B1 => n8882, B2 => 
                           n9662, ZN => n3378);
   U2514 : OAI22_X1 port map( A1 => n9269, A2 => n9659, B1 => n8883, B2 => 
                           n9662, ZN => n3379);
   U2515 : OAI22_X1 port map( A1 => n9266, A2 => n9659, B1 => n8884, B2 => 
                           n9662, ZN => n3380);
   U2516 : OAI22_X1 port map( A1 => n9263, A2 => n9659, B1 => n8885, B2 => 
                           n9662, ZN => n3381);
   U2517 : OAI22_X1 port map( A1 => n9260, A2 => n9592, B1 => n8295, B2 => 
                           n9595, ZN => n3190);
   U2518 : OAI22_X1 port map( A1 => n9257, A2 => n9593, B1 => n8296, B2 => 
                           n9595, ZN => n3191);
   U2519 : OAI22_X1 port map( A1 => n9254, A2 => n9592, B1 => n8297, B2 => 
                           n9595, ZN => n3192);
   U2520 : OAI22_X1 port map( A1 => n9251, A2 => n9593, B1 => n8298, B2 => 
                           n9595, ZN => n3193);
   U2521 : OAI22_X1 port map( A1 => n9248, A2 => n9592, B1 => n8299, B2 => 
                           n9594, ZN => n3194);
   U2522 : OAI22_X1 port map( A1 => n9245, A2 => n9593, B1 => n8300, B2 => 
                           n9594, ZN => n3195);
   U2523 : OAI22_X1 port map( A1 => n9242, A2 => n9592, B1 => n8301, B2 => 
                           n9594, ZN => n3196);
   U2524 : OAI22_X1 port map( A1 => n9239, A2 => n9593, B1 => n8302, B2 => 
                           n9594, ZN => n3197);
   U2525 : OAI22_X1 port map( A1 => n9329, A2 => n9592, B1 => n8631, B2 => 
                           n9601, ZN => n3167);
   U2526 : OAI22_X1 port map( A1 => n9326, A2 => n9592, B1 => n8632, B2 => 
                           n9601, ZN => n3168);
   U2527 : OAI22_X1 port map( A1 => n9323, A2 => n9592, B1 => n8633, B2 => 
                           n9601, ZN => n3169);
   U2528 : OAI22_X1 port map( A1 => n9320, A2 => n9592, B1 => n8634, B2 => 
                           n9600, ZN => n3170);
   U2529 : OAI22_X1 port map( A1 => n9317, A2 => n9592, B1 => n8635, B2 => 
                           n9600, ZN => n3171);
   U2530 : OAI22_X1 port map( A1 => n9311, A2 => n9592, B1 => n8637, B2 => 
                           n9600, ZN => n3173);
   U2531 : OAI22_X1 port map( A1 => n9308, A2 => n9592, B1 => n8638, B2 => 
                           n9599, ZN => n3174);
   U2532 : OAI22_X1 port map( A1 => n9305, A2 => n9592, B1 => n8639, B2 => 
                           n9599, ZN => n3175);
   U2533 : OAI22_X1 port map( A1 => n9302, A2 => n9592, B1 => n8640, B2 => 
                           n9599, ZN => n3176);
   U2534 : OAI22_X1 port map( A1 => n9299, A2 => n9592, B1 => n8641, B2 => 
                           n9599, ZN => n3177);
   U2535 : OAI22_X1 port map( A1 => n9296, A2 => n9593, B1 => n8642, B2 => 
                           n9598, ZN => n3178);
   U2536 : OAI22_X1 port map( A1 => n9290, A2 => n9593, B1 => n8644, B2 => 
                           n9598, ZN => n3180);
   U2537 : OAI22_X1 port map( A1 => n9287, A2 => n9593, B1 => n8645, B2 => 
                           n9598, ZN => n3181);
   U2538 : OAI22_X1 port map( A1 => n9284, A2 => n9593, B1 => n8646, B2 => 
                           n9597, ZN => n3182);
   U2539 : OAI22_X1 port map( A1 => n9278, A2 => n9593, B1 => n8648, B2 => 
                           n9597, ZN => n3184);
   U2540 : OAI22_X1 port map( A1 => n9275, A2 => n9593, B1 => n8649, B2 => 
                           n9597, ZN => n3185);
   U2541 : OAI22_X1 port map( A1 => n9272, A2 => n9593, B1 => n8650, B2 => 
                           n9596, ZN => n3186);
   U2542 : OAI22_X1 port map( A1 => n9269, A2 => n9593, B1 => n8651, B2 => 
                           n9596, ZN => n3187);
   U2543 : OAI22_X1 port map( A1 => n9266, A2 => n9593, B1 => n8652, B2 => 
                           n9596, ZN => n3188);
   U2544 : OAI22_X1 port map( A1 => n9263, A2 => n9593, B1 => n8653, B2 => 
                           n9596, ZN => n3189);
   U2545 : OAI22_X1 port map( A1 => n9332, A2 => n9603, B1 => n8654, B2 => 
                           n9612, ZN => n3198);
   U2546 : OAI22_X1 port map( A1 => n9314, A2 => n9603, B1 => n8660, B2 => 
                           n9611, ZN => n3204);
   U2547 : OAI22_X1 port map( A1 => n9293, A2 => n9604, B1 => n8667, B2 => 
                           n9609, ZN => n3211);
   U2548 : OAI22_X1 port map( A1 => n9281, A2 => n9604, B1 => n8671, B2 => 
                           n9608, ZN => n3215);
   U2549 : OAI22_X1 port map( A1 => n9333, A2 => n9581, B1 => n8566, B2 => 
                           n9590, ZN => n3134);
   U2550 : OAI22_X1 port map( A1 => n9332, A2 => n9724, B1 => n8598, B2 => 
                           n9726, ZN => n3952);
   U2551 : OAI22_X1 port map( A1 => n9331, A2 => n9812, B1 => n8245, B2 => 
                           n9821, ZN => n9014);
   U2552 : OAI22_X1 port map( A1 => n9313, A2 => n9812, B1 => n8233, B2 => 
                           n9820, ZN => n9020);
   U2553 : OAI22_X1 port map( A1 => n9292, A2 => n9813, B1 => n8219, B2 => 
                           n9818, ZN => n9027);
   U2554 : OAI22_X1 port map( A1 => n9280, A2 => n9813, B1 => n8211, B2 => 
                           n9817, ZN => n9031);
   U2555 : OAI22_X1 port map( A1 => n9332, A2 => n9636, B1 => n8774, B2 => 
                           n9645, ZN => n3294);
   U2556 : OAI22_X1 port map( A1 => n9314, A2 => n9636, B1 => n8780, B2 => 
                           n9644, ZN => n3300);
   U2557 : OAI22_X1 port map( A1 => n9293, A2 => n9637, B1 => n8787, B2 => 
                           n9642, ZN => n3307);
   U2558 : OAI22_X1 port map( A1 => n9281, A2 => n9637, B1 => n8791, B2 => 
                           n9641, ZN => n3311);
   U2559 : OAI22_X1 port map( A1 => n9332, A2 => n9592, B1 => n8630, B2 => 
                           n9601, ZN => n3166);
   U2560 : OAI22_X1 port map( A1 => n9314, A2 => n9592, B1 => n8636, B2 => 
                           n9600, ZN => n3172);
   U2561 : OAI22_X1 port map( A1 => n9293, A2 => n9593, B1 => n8643, B2 => 
                           n9598, ZN => n3179);
   U2562 : OAI22_X1 port map( A1 => n9281, A2 => n9593, B1 => n8647, B2 => 
                           n9597, ZN => n3183);
   U2563 : OAI22_X1 port map( A1 => n9333, A2 => n9526, B1 => n8263, B2 => 
                           n9535, ZN => n2942);
   U2564 : OAI22_X1 port map( A1 => n9330, A2 => n9526, B1 => n8264, B2 => 
                           n9535, ZN => n2943);
   U2565 : OAI22_X1 port map( A1 => n9327, A2 => n9526, B1 => n8265, B2 => 
                           n9535, ZN => n2944);
   U2566 : OAI22_X1 port map( A1 => n9324, A2 => n9526, B1 => n8266, B2 => 
                           n9535, ZN => n2945);
   U2567 : OAI22_X1 port map( A1 => n9321, A2 => n9526, B1 => n8267, B2 => 
                           n9534, ZN => n2946);
   U2568 : OAI22_X1 port map( A1 => n9318, A2 => n9526, B1 => n8268, B2 => 
                           n9534, ZN => n2947);
   U2569 : OAI22_X1 port map( A1 => n9315, A2 => n9526, B1 => n8269, B2 => 
                           n9534, ZN => n2948);
   U2570 : OAI22_X1 port map( A1 => n9312, A2 => n9526, B1 => n8270, B2 => 
                           n9534, ZN => n2949);
   U2571 : OAI22_X1 port map( A1 => n9309, A2 => n9526, B1 => n8271, B2 => 
                           n9533, ZN => n2950);
   U2572 : OAI22_X1 port map( A1 => n9306, A2 => n9526, B1 => n8272, B2 => 
                           n9533, ZN => n2951);
   U2573 : OAI22_X1 port map( A1 => n9303, A2 => n9526, B1 => n8273, B2 => 
                           n9533, ZN => n2952);
   U2574 : OAI22_X1 port map( A1 => n9300, A2 => n9526, B1 => n8274, B2 => 
                           n9533, ZN => n2953);
   U2575 : OAI22_X1 port map( A1 => n9297, A2 => n9527, B1 => n8275, B2 => 
                           n9532, ZN => n2954);
   U2576 : OAI22_X1 port map( A1 => n9294, A2 => n9527, B1 => n8276, B2 => 
                           n9532, ZN => n2955);
   U2577 : OAI22_X1 port map( A1 => n9291, A2 => n9527, B1 => n8277, B2 => 
                           n9532, ZN => n2956);
   U2578 : OAI22_X1 port map( A1 => n9288, A2 => n9527, B1 => n8278, B2 => 
                           n9532, ZN => n2957);
   U2579 : OAI22_X1 port map( A1 => n9285, A2 => n9527, B1 => n8279, B2 => 
                           n9531, ZN => n2958);
   U2580 : OAI22_X1 port map( A1 => n9282, A2 => n9527, B1 => n8280, B2 => 
                           n9531, ZN => n2959);
   U2581 : OAI22_X1 port map( A1 => n9279, A2 => n9527, B1 => n8281, B2 => 
                           n9531, ZN => n2960);
   U2582 : OAI22_X1 port map( A1 => n9276, A2 => n9527, B1 => n8282, B2 => 
                           n9531, ZN => n2961);
   U2583 : OAI22_X1 port map( A1 => n9273, A2 => n9527, B1 => n8283, B2 => 
                           n9530, ZN => n2962);
   U2584 : OAI22_X1 port map( A1 => n9270, A2 => n9527, B1 => n8284, B2 => 
                           n9530, ZN => n2963);
   U2585 : OAI22_X1 port map( A1 => n9267, A2 => n9527, B1 => n8285, B2 => 
                           n9530, ZN => n2964);
   U2586 : OAI22_X1 port map( A1 => n9264, A2 => n9527, B1 => n8286, B2 => 
                           n9530, ZN => n2965);
   U2587 : OAI22_X1 port map( A1 => n9333, A2 => n9537, B1 => n2350, B2 => 
                           n9546, ZN => n2974);
   U2588 : OAI22_X1 port map( A1 => n9330, A2 => n9537, B1 => n2342, B2 => 
                           n9546, ZN => n2975);
   U2589 : OAI22_X1 port map( A1 => n9327, A2 => n9537, B1 => n2334, B2 => 
                           n9546, ZN => n2976);
   U2590 : OAI22_X1 port map( A1 => n9324, A2 => n9537, B1 => n2326, B2 => 
                           n9546, ZN => n2977);
   U2591 : OAI22_X1 port map( A1 => n9321, A2 => n9537, B1 => n2318, B2 => 
                           n9545, ZN => n2978);
   U2592 : OAI22_X1 port map( A1 => n9318, A2 => n9537, B1 => n2310, B2 => 
                           n9545, ZN => n2979);
   U2593 : OAI22_X1 port map( A1 => n9315, A2 => n9537, B1 => n2302, B2 => 
                           n9545, ZN => n2980);
   U2594 : OAI22_X1 port map( A1 => n9312, A2 => n9537, B1 => n2294, B2 => 
                           n9545, ZN => n2981);
   U2595 : OAI22_X1 port map( A1 => n9309, A2 => n9537, B1 => n2286, B2 => 
                           n9544, ZN => n2982);
   U2596 : OAI22_X1 port map( A1 => n9306, A2 => n9537, B1 => n2278, B2 => 
                           n9544, ZN => n2983);
   U2597 : OAI22_X1 port map( A1 => n9303, A2 => n9537, B1 => n2270, B2 => 
                           n9544, ZN => n2984);
   U2598 : OAI22_X1 port map( A1 => n9300, A2 => n9537, B1 => n2262, B2 => 
                           n9544, ZN => n2985);
   U2599 : OAI22_X1 port map( A1 => n9297, A2 => n9538, B1 => n2254, B2 => 
                           n9543, ZN => n2986);
   U2600 : OAI22_X1 port map( A1 => n9294, A2 => n9538, B1 => n2246, B2 => 
                           n9543, ZN => n2987);
   U2601 : OAI22_X1 port map( A1 => n9291, A2 => n9538, B1 => n2238, B2 => 
                           n9543, ZN => n2988);
   U2602 : OAI22_X1 port map( A1 => n9288, A2 => n9538, B1 => n2230, B2 => 
                           n9543, ZN => n2989);
   U2603 : OAI22_X1 port map( A1 => n9285, A2 => n9538, B1 => n2222, B2 => 
                           n9542, ZN => n2990);
   U2604 : OAI22_X1 port map( A1 => n9282, A2 => n9538, B1 => n2214, B2 => 
                           n9542, ZN => n2991);
   U2605 : OAI22_X1 port map( A1 => n9279, A2 => n9538, B1 => n2206, B2 => 
                           n9542, ZN => n2992);
   U2606 : OAI22_X1 port map( A1 => n9276, A2 => n9538, B1 => n2198, B2 => 
                           n9542, ZN => n2993);
   U2607 : OAI22_X1 port map( A1 => n9273, A2 => n9538, B1 => n2190, B2 => 
                           n9541, ZN => n2994);
   U2608 : OAI22_X1 port map( A1 => n9270, A2 => n9538, B1 => n2182, B2 => 
                           n9541, ZN => n2995);
   U2609 : OAI22_X1 port map( A1 => n9267, A2 => n9538, B1 => n2174, B2 => 
                           n9541, ZN => n2996);
   U2610 : OAI22_X1 port map( A1 => n9264, A2 => n9538, B1 => n2166, B2 => 
                           n9541, ZN => n2997);
   U2611 : OAI22_X1 port map( A1 => n9261, A2 => n9526, B1 => n8335, B2 => 
                           n9529, ZN => n2966);
   U2612 : OAI22_X1 port map( A1 => n9258, A2 => n9527, B1 => n8336, B2 => 
                           n9529, ZN => n2967);
   U2613 : OAI22_X1 port map( A1 => n9255, A2 => n9526, B1 => n8337, B2 => 
                           n9529, ZN => n2968);
   U2614 : OAI22_X1 port map( A1 => n9252, A2 => n9527, B1 => n8338, B2 => 
                           n9529, ZN => n2969);
   U2615 : OAI22_X1 port map( A1 => n9249, A2 => n9526, B1 => n8339, B2 => 
                           n9528, ZN => n2970);
   U2616 : OAI22_X1 port map( A1 => n9246, A2 => n9527, B1 => n8340, B2 => 
                           n9528, ZN => n2971);
   U2617 : OAI22_X1 port map( A1 => n9243, A2 => n9526, B1 => n8341, B2 => 
                           n9528, ZN => n2972);
   U2618 : OAI22_X1 port map( A1 => n9240, A2 => n9527, B1 => n8342, B2 => 
                           n9528, ZN => n2973);
   U2619 : OAI22_X1 port map( A1 => n9261, A2 => n9537, B1 => n2158, B2 => 
                           n9540, ZN => n2998);
   U2620 : OAI22_X1 port map( A1 => n9258, A2 => n9538, B1 => n2150, B2 => 
                           n9540, ZN => n2999);
   U2621 : OAI22_X1 port map( A1 => n9255, A2 => n9537, B1 => n2142, B2 => 
                           n9540, ZN => n3000);
   U2622 : OAI22_X1 port map( A1 => n9252, A2 => n9538, B1 => n2134, B2 => 
                           n9540, ZN => n3001);
   U2623 : OAI22_X1 port map( A1 => n9249, A2 => n9537, B1 => n2126, B2 => 
                           n9539, ZN => n3002);
   U2624 : OAI22_X1 port map( A1 => n9246, A2 => n9538, B1 => n2118, B2 => 
                           n9539, ZN => n3003);
   U2625 : OAI22_X1 port map( A1 => n9243, A2 => n9537, B1 => n2110, B2 => 
                           n9539, ZN => n3004);
   U2626 : OAI22_X1 port map( A1 => n9240, A2 => n9538, B1 => n2102, B2 => 
                           n9539, ZN => n3005);
   U2627 : OAI22_X1 port map( A1 => n9331, A2 => n9856, B1 => n2348, B2 => 
                           n9865, ZN => n9142);
   U2628 : OAI22_X1 port map( A1 => n9328, A2 => n9856, B1 => n2340, B2 => 
                           n9865, ZN => n9143);
   U2629 : OAI22_X1 port map( A1 => n9325, A2 => n9856, B1 => n2332, B2 => 
                           n9865, ZN => n9144);
   U2630 : OAI22_X1 port map( A1 => n9322, A2 => n9856, B1 => n2324, B2 => 
                           n9865, ZN => n9145);
   U2631 : OAI22_X1 port map( A1 => n9319, A2 => n9856, B1 => n2316, B2 => 
                           n9864, ZN => n9146);
   U2632 : OAI22_X1 port map( A1 => n9316, A2 => n9856, B1 => n2308, B2 => 
                           n9864, ZN => n9147);
   U2633 : OAI22_X1 port map( A1 => n9313, A2 => n9856, B1 => n2300, B2 => 
                           n9864, ZN => n9148);
   U2634 : OAI22_X1 port map( A1 => n9310, A2 => n9856, B1 => n2292, B2 => 
                           n9864, ZN => n9149);
   U2635 : OAI22_X1 port map( A1 => n9307, A2 => n9856, B1 => n2284, B2 => 
                           n9863, ZN => n9150);
   U2636 : OAI22_X1 port map( A1 => n9304, A2 => n9856, B1 => n2276, B2 => 
                           n9863, ZN => n9151);
   U2637 : OAI22_X1 port map( A1 => n9301, A2 => n9856, B1 => n2268, B2 => 
                           n9863, ZN => n9152);
   U2638 : OAI22_X1 port map( A1 => n9298, A2 => n9856, B1 => n2260, B2 => 
                           n9863, ZN => n9153);
   U2639 : OAI22_X1 port map( A1 => n9295, A2 => n9857, B1 => n2252, B2 => 
                           n9862, ZN => n9154);
   U2640 : OAI22_X1 port map( A1 => n9292, A2 => n9857, B1 => n2244, B2 => 
                           n9862, ZN => n9155);
   U2641 : OAI22_X1 port map( A1 => n9289, A2 => n9857, B1 => n2236, B2 => 
                           n9862, ZN => n9156);
   U2642 : OAI22_X1 port map( A1 => n9286, A2 => n9857, B1 => n2228, B2 => 
                           n9862, ZN => n9157);
   U2643 : OAI22_X1 port map( A1 => n9283, A2 => n9857, B1 => n2220, B2 => 
                           n9861, ZN => n9158);
   U2644 : OAI22_X1 port map( A1 => n9280, A2 => n9857, B1 => n2212, B2 => 
                           n9861, ZN => n9159);
   U2645 : OAI22_X1 port map( A1 => n9277, A2 => n9857, B1 => n2204, B2 => 
                           n9861, ZN => n9160);
   U2646 : OAI22_X1 port map( A1 => n9274, A2 => n9857, B1 => n2196, B2 => 
                           n9861, ZN => n9161);
   U2647 : OAI22_X1 port map( A1 => n9271, A2 => n9857, B1 => n2188, B2 => 
                           n9860, ZN => n9162);
   U2648 : OAI22_X1 port map( A1 => n9268, A2 => n9857, B1 => n2180, B2 => 
                           n9860, ZN => n9163);
   U2649 : OAI22_X1 port map( A1 => n9265, A2 => n9857, B1 => n2172, B2 => 
                           n9860, ZN => n9164);
   U2650 : OAI22_X1 port map( A1 => n9262, A2 => n9857, B1 => n2164, B2 => 
                           n9860, ZN => n9165);
   U2651 : OAI22_X1 port map( A1 => n9259, A2 => n9856, B1 => n2156, B2 => 
                           n9859, ZN => n9166);
   U2652 : OAI22_X1 port map( A1 => n9256, A2 => n9857, B1 => n2148, B2 => 
                           n9859, ZN => n9167);
   U2653 : OAI22_X1 port map( A1 => n9253, A2 => n9856, B1 => n2140, B2 => 
                           n9859, ZN => n9168);
   U2654 : OAI22_X1 port map( A1 => n9250, A2 => n9857, B1 => n2132, B2 => 
                           n9859, ZN => n9169);
   U2655 : OAI22_X1 port map( A1 => n9247, A2 => n9856, B1 => n2124, B2 => 
                           n9858, ZN => n9170);
   U2656 : OAI22_X1 port map( A1 => n9244, A2 => n9857, B1 => n2116, B2 => 
                           n9858, ZN => n9171);
   U2657 : OAI22_X1 port map( A1 => n9241, A2 => n9856, B1 => n2108, B2 => 
                           n9858, ZN => n9172);
   U2658 : OAI22_X1 port map( A1 => n9238, A2 => n9857, B1 => n2100, B2 => 
                           n9858, ZN => n9173);
   U2659 : OAI22_X1 port map( A1 => n9331, A2 => n9823, B1 => n2355, B2 => 
                           n9832, ZN => n9046);
   U2660 : OAI22_X1 port map( A1 => n9328, A2 => n9823, B1 => n2347, B2 => 
                           n9832, ZN => n9047);
   U2661 : OAI22_X1 port map( A1 => n9325, A2 => n9823, B1 => n2339, B2 => 
                           n9832, ZN => n9048);
   U2662 : OAI22_X1 port map( A1 => n9322, A2 => n9823, B1 => n2331, B2 => 
                           n9832, ZN => n9049);
   U2663 : OAI22_X1 port map( A1 => n9319, A2 => n9823, B1 => n2323, B2 => 
                           n9831, ZN => n9050);
   U2664 : OAI22_X1 port map( A1 => n9316, A2 => n9823, B1 => n2315, B2 => 
                           n9831, ZN => n9051);
   U2665 : OAI22_X1 port map( A1 => n9313, A2 => n9823, B1 => n2307, B2 => 
                           n9831, ZN => n9052);
   U2666 : OAI22_X1 port map( A1 => n9310, A2 => n9823, B1 => n2299, B2 => 
                           n9831, ZN => n9053);
   U2667 : OAI22_X1 port map( A1 => n9307, A2 => n9823, B1 => n2291, B2 => 
                           n9830, ZN => n9054);
   U2668 : OAI22_X1 port map( A1 => n9304, A2 => n9823, B1 => n2283, B2 => 
                           n9830, ZN => n9055);
   U2669 : OAI22_X1 port map( A1 => n9301, A2 => n9823, B1 => n2275, B2 => 
                           n9830, ZN => n9056);
   U2670 : OAI22_X1 port map( A1 => n9298, A2 => n9823, B1 => n2267, B2 => 
                           n9830, ZN => n9057);
   U2671 : OAI22_X1 port map( A1 => n9295, A2 => n9824, B1 => n2259, B2 => 
                           n9829, ZN => n9058);
   U2672 : OAI22_X1 port map( A1 => n9292, A2 => n9824, B1 => n2251, B2 => 
                           n9829, ZN => n9059);
   U2673 : OAI22_X1 port map( A1 => n9289, A2 => n9824, B1 => n2243, B2 => 
                           n9829, ZN => n9060);
   U2674 : OAI22_X1 port map( A1 => n9286, A2 => n9824, B1 => n2235, B2 => 
                           n9829, ZN => n9061);
   U2675 : OAI22_X1 port map( A1 => n9283, A2 => n9824, B1 => n2227, B2 => 
                           n9828, ZN => n9062);
   U2676 : OAI22_X1 port map( A1 => n9280, A2 => n9824, B1 => n2219, B2 => 
                           n9828, ZN => n9063);
   U2677 : OAI22_X1 port map( A1 => n9277, A2 => n9824, B1 => n2211, B2 => 
                           n9828, ZN => n9064);
   U2678 : OAI22_X1 port map( A1 => n9274, A2 => n9824, B1 => n2203, B2 => 
                           n9828, ZN => n9065);
   U2679 : OAI22_X1 port map( A1 => n9271, A2 => n9824, B1 => n2195, B2 => 
                           n9827, ZN => n9066);
   U2680 : OAI22_X1 port map( A1 => n9268, A2 => n9824, B1 => n2187, B2 => 
                           n9827, ZN => n9067);
   U2681 : OAI22_X1 port map( A1 => n9265, A2 => n9824, B1 => n2179, B2 => 
                           n9827, ZN => n9068);
   U2682 : OAI22_X1 port map( A1 => n9262, A2 => n9824, B1 => n2171, B2 => 
                           n9827, ZN => n9069);
   U2683 : OAI22_X1 port map( A1 => n9259, A2 => n9823, B1 => n2163, B2 => 
                           n9826, ZN => n9070);
   U2684 : OAI22_X1 port map( A1 => n9256, A2 => n9824, B1 => n2155, B2 => 
                           n9826, ZN => n9071);
   U2685 : OAI22_X1 port map( A1 => n9253, A2 => n9823, B1 => n2147, B2 => 
                           n9826, ZN => n9072);
   U2686 : OAI22_X1 port map( A1 => n9250, A2 => n9824, B1 => n2139, B2 => 
                           n9826, ZN => n9073);
   U2687 : OAI22_X1 port map( A1 => n9247, A2 => n9823, B1 => n2131, B2 => 
                           n9825, ZN => n9074);
   U2688 : OAI22_X1 port map( A1 => n9244, A2 => n9824, B1 => n2123, B2 => 
                           n9825, ZN => n9075);
   U2689 : OAI22_X1 port map( A1 => n9241, A2 => n9823, B1 => n2115, B2 => 
                           n9825, ZN => n9076);
   U2690 : OAI22_X1 port map( A1 => n9238, A2 => n9824, B1 => n2107, B2 => 
                           n9825, ZN => n9077);
   U2691 : OAI22_X1 port map( A1 => n9332, A2 => n9714, B1 => n8686, B2 => 
                           n9715, ZN => n3949);
   U2692 : OAI22_X1 port map( A1 => n9329, A2 => n9713, B1 => n8687, B2 => 
                           n9715, ZN => n3933);
   U2693 : OAI22_X1 port map( A1 => n9326, A2 => n9714, B1 => n8688, B2 => 
                           n9715, ZN => n3917);
   U2694 : OAI22_X1 port map( A1 => n9323, A2 => n9713, B1 => n8689, B2 => 
                           n9715, ZN => n3901);
   U2695 : OAI22_X1 port map( A1 => n9320, A2 => n9714, B1 => n8690, B2 => 
                           n9716, ZN => n3885);
   U2696 : OAI22_X1 port map( A1 => n9317, A2 => n9713, B1 => n8691, B2 => 
                           n9716, ZN => n3869);
   U2697 : OAI22_X1 port map( A1 => n9314, A2 => n9714, B1 => n8692, B2 => 
                           n9716, ZN => n3853);
   U2698 : OAI22_X1 port map( A1 => n9311, A2 => n9713, B1 => n8693, B2 => 
                           n9716, ZN => n3837);
   U2699 : OAI22_X1 port map( A1 => n9308, A2 => n9714, B1 => n8694, B2 => 
                           n9717, ZN => n3821);
   U2700 : OAI22_X1 port map( A1 => n9305, A2 => n9714, B1 => n8695, B2 => 
                           n9717, ZN => n3805);
   U2701 : OAI22_X1 port map( A1 => n9302, A2 => n9714, B1 => n8696, B2 => 
                           n9717, ZN => n3789);
   U2702 : OAI22_X1 port map( A1 => n9299, A2 => n9714, B1 => n8697, B2 => 
                           n9717, ZN => n3773);
   U2703 : OAI22_X1 port map( A1 => n9296, A2 => n9714, B1 => n8698, B2 => 
                           n9718, ZN => n3757);
   U2704 : OAI22_X1 port map( A1 => n9293, A2 => n9714, B1 => n8699, B2 => 
                           n9718, ZN => n3741);
   U2705 : OAI22_X1 port map( A1 => n9290, A2 => n9714, B1 => n8700, B2 => 
                           n9718, ZN => n3725);
   U2706 : OAI22_X1 port map( A1 => n9287, A2 => n9714, B1 => n8701, B2 => 
                           n9718, ZN => n3709);
   U2707 : OAI22_X1 port map( A1 => n9284, A2 => n9714, B1 => n8702, B2 => 
                           n9719, ZN => n3693);
   U2708 : OAI22_X1 port map( A1 => n9281, A2 => n9714, B1 => n8703, B2 => 
                           n9719, ZN => n3677);
   U2709 : OAI22_X1 port map( A1 => n9278, A2 => n9714, B1 => n8704, B2 => 
                           n9719, ZN => n3661);
   U2710 : OAI22_X1 port map( A1 => n9275, A2 => n9714, B1 => n8705, B2 => 
                           n9719, ZN => n3645);
   U2711 : OAI22_X1 port map( A1 => n9272, A2 => n9713, B1 => n8706, B2 => 
                           n9720, ZN => n3629);
   U2712 : OAI22_X1 port map( A1 => n9269, A2 => n9713, B1 => n8707, B2 => 
                           n9720, ZN => n3613);
   U2713 : OAI22_X1 port map( A1 => n9266, A2 => n9713, B1 => n8708, B2 => 
                           n9720, ZN => n3597);
   U2714 : OAI22_X1 port map( A1 => n9263, A2 => n9713, B1 => n8709, B2 => 
                           n9720, ZN => n3581);
   U2715 : OAI22_X1 port map( A1 => n9260, A2 => n9713, B1 => n8710, B2 => 
                           n9721, ZN => n3565);
   U2716 : OAI22_X1 port map( A1 => n9257, A2 => n9713, B1 => n8711, B2 => 
                           n9721, ZN => n3549);
   U2717 : OAI22_X1 port map( A1 => n9254, A2 => n9713, B1 => n8712, B2 => 
                           n9721, ZN => n3533);
   U2718 : OAI22_X1 port map( A1 => n9251, A2 => n9713, B1 => n8713, B2 => 
                           n9721, ZN => n3517);
   U2719 : OAI22_X1 port map( A1 => n9248, A2 => n9713, B1 => n8714, B2 => 
                           n9722, ZN => n3501);
   U2720 : OAI22_X1 port map( A1 => n9245, A2 => n9713, B1 => n8715, B2 => 
                           n9722, ZN => n3485);
   U2721 : OAI22_X1 port map( A1 => n9242, A2 => n9713, B1 => n8716, B2 => 
                           n9722, ZN => n3469);
   U2722 : OAI22_X1 port map( A1 => n9239, A2 => n9713, B1 => n8717, B2 => 
                           n9722, ZN => n3453);
   U2723 : OAI22_X1 port map( A1 => n9332, A2 => n9703, B1 => n2354, B2 => 
                           n9704, ZN => n3948);
   U2724 : OAI22_X1 port map( A1 => n9329, A2 => n9702, B1 => n2346, B2 => 
                           n9704, ZN => n3932);
   U2725 : OAI22_X1 port map( A1 => n9326, A2 => n9703, B1 => n2338, B2 => 
                           n9704, ZN => n3916);
   U2726 : OAI22_X1 port map( A1 => n9323, A2 => n9702, B1 => n2330, B2 => 
                           n9704, ZN => n3900);
   U2727 : OAI22_X1 port map( A1 => n9320, A2 => n9703, B1 => n2322, B2 => 
                           n9705, ZN => n3884);
   U2728 : OAI22_X1 port map( A1 => n9317, A2 => n9702, B1 => n2314, B2 => 
                           n9705, ZN => n3868);
   U2729 : OAI22_X1 port map( A1 => n9314, A2 => n9703, B1 => n2306, B2 => 
                           n9705, ZN => n3852);
   U2730 : OAI22_X1 port map( A1 => n9311, A2 => n9702, B1 => n2298, B2 => 
                           n9705, ZN => n3836);
   U2731 : OAI22_X1 port map( A1 => n9308, A2 => n9703, B1 => n2290, B2 => 
                           n9706, ZN => n3820);
   U2732 : OAI22_X1 port map( A1 => n9305, A2 => n9703, B1 => n2282, B2 => 
                           n9706, ZN => n3804);
   U2733 : OAI22_X1 port map( A1 => n9302, A2 => n9703, B1 => n2274, B2 => 
                           n9706, ZN => n3788);
   U2734 : OAI22_X1 port map( A1 => n9299, A2 => n9703, B1 => n2266, B2 => 
                           n9706, ZN => n3772);
   U2735 : OAI22_X1 port map( A1 => n9296, A2 => n9703, B1 => n2258, B2 => 
                           n9707, ZN => n3756);
   U2736 : OAI22_X1 port map( A1 => n9293, A2 => n9703, B1 => n2250, B2 => 
                           n9707, ZN => n3740);
   U2737 : OAI22_X1 port map( A1 => n9290, A2 => n9703, B1 => n2242, B2 => 
                           n9707, ZN => n3724);
   U2738 : OAI22_X1 port map( A1 => n9287, A2 => n9703, B1 => n2234, B2 => 
                           n9707, ZN => n3708);
   U2739 : OAI22_X1 port map( A1 => n9284, A2 => n9703, B1 => n2226, B2 => 
                           n9708, ZN => n3692);
   U2740 : OAI22_X1 port map( A1 => n9281, A2 => n9703, B1 => n2218, B2 => 
                           n9708, ZN => n3676);
   U2741 : OAI22_X1 port map( A1 => n9278, A2 => n9703, B1 => n2210, B2 => 
                           n9708, ZN => n3660);
   U2742 : OAI22_X1 port map( A1 => n9275, A2 => n9703, B1 => n2202, B2 => 
                           n9708, ZN => n3644);
   U2743 : OAI22_X1 port map( A1 => n9272, A2 => n9702, B1 => n2194, B2 => 
                           n9709, ZN => n3628);
   U2744 : OAI22_X1 port map( A1 => n9269, A2 => n9702, B1 => n2186, B2 => 
                           n9709, ZN => n3612);
   U2745 : OAI22_X1 port map( A1 => n9266, A2 => n9702, B1 => n2178, B2 => 
                           n9709, ZN => n3596);
   U2746 : OAI22_X1 port map( A1 => n9263, A2 => n9702, B1 => n2170, B2 => 
                           n9709, ZN => n3580);
   U2747 : OAI22_X1 port map( A1 => n9260, A2 => n9702, B1 => n2162, B2 => 
                           n9710, ZN => n3564);
   U2748 : OAI22_X1 port map( A1 => n9257, A2 => n9702, B1 => n2154, B2 => 
                           n9710, ZN => n3548);
   U2749 : OAI22_X1 port map( A1 => n9254, A2 => n9702, B1 => n2146, B2 => 
                           n9710, ZN => n3532);
   U2750 : OAI22_X1 port map( A1 => n9251, A2 => n9702, B1 => n2138, B2 => 
                           n9710, ZN => n3516);
   U2751 : OAI22_X1 port map( A1 => n9248, A2 => n9702, B1 => n2130, B2 => 
                           n9711, ZN => n3500);
   U2752 : OAI22_X1 port map( A1 => n9245, A2 => n9702, B1 => n2122, B2 => 
                           n9711, ZN => n3484);
   U2753 : OAI22_X1 port map( A1 => n9242, A2 => n9702, B1 => n2114, B2 => 
                           n9711, ZN => n3468);
   U2754 : OAI22_X1 port map( A1 => n9239, A2 => n9702, B1 => n2106, B2 => 
                           n9711, ZN => n3452);
   U2755 : OAI22_X1 port map( A1 => n9331, A2 => n9801, B1 => n2353, B2 => 
                           n9810, ZN => n8982);
   U2756 : OAI22_X1 port map( A1 => n9328, A2 => n9801, B1 => n2345, B2 => 
                           n9810, ZN => n8983);
   U2757 : OAI22_X1 port map( A1 => n9325, A2 => n9801, B1 => n2337, B2 => 
                           n9810, ZN => n8984);
   U2758 : OAI22_X1 port map( A1 => n9322, A2 => n9801, B1 => n2329, B2 => 
                           n9810, ZN => n8985);
   U2759 : OAI22_X1 port map( A1 => n9319, A2 => n9801, B1 => n2321, B2 => 
                           n9809, ZN => n8986);
   U2760 : OAI22_X1 port map( A1 => n9316, A2 => n9801, B1 => n2313, B2 => 
                           n9809, ZN => n8987);
   U2761 : OAI22_X1 port map( A1 => n9313, A2 => n9801, B1 => n2305, B2 => 
                           n9809, ZN => n8988);
   U2762 : OAI22_X1 port map( A1 => n9310, A2 => n9801, B1 => n2297, B2 => 
                           n9809, ZN => n8989);
   U2763 : OAI22_X1 port map( A1 => n9307, A2 => n9801, B1 => n2289, B2 => 
                           n9808, ZN => n8990);
   U2764 : OAI22_X1 port map( A1 => n9304, A2 => n9801, B1 => n2281, B2 => 
                           n9808, ZN => n8991);
   U2765 : OAI22_X1 port map( A1 => n9301, A2 => n9801, B1 => n2273, B2 => 
                           n9808, ZN => n8992);
   U2766 : OAI22_X1 port map( A1 => n9298, A2 => n9801, B1 => n2265, B2 => 
                           n9808, ZN => n8993);
   U2767 : OAI22_X1 port map( A1 => n9295, A2 => n9802, B1 => n2257, B2 => 
                           n9807, ZN => n8994);
   U2768 : OAI22_X1 port map( A1 => n9292, A2 => n9802, B1 => n2249, B2 => 
                           n9807, ZN => n8995);
   U2769 : OAI22_X1 port map( A1 => n9289, A2 => n9802, B1 => n2241, B2 => 
                           n9807, ZN => n8996);
   U2770 : OAI22_X1 port map( A1 => n9286, A2 => n9802, B1 => n2233, B2 => 
                           n9807, ZN => n8997);
   U2771 : OAI22_X1 port map( A1 => n9283, A2 => n9802, B1 => n2225, B2 => 
                           n9806, ZN => n8998);
   U2772 : OAI22_X1 port map( A1 => n9280, A2 => n9802, B1 => n2217, B2 => 
                           n9806, ZN => n8999);
   U2773 : OAI22_X1 port map( A1 => n9277, A2 => n9802, B1 => n2209, B2 => 
                           n9806, ZN => n9000);
   U2774 : OAI22_X1 port map( A1 => n9274, A2 => n9802, B1 => n2201, B2 => 
                           n9806, ZN => n9001);
   U2775 : OAI22_X1 port map( A1 => n9271, A2 => n9802, B1 => n2193, B2 => 
                           n9805, ZN => n9002);
   U2776 : OAI22_X1 port map( A1 => n9268, A2 => n9802, B1 => n2185, B2 => 
                           n9805, ZN => n9003);
   U2777 : OAI22_X1 port map( A1 => n9265, A2 => n9802, B1 => n2177, B2 => 
                           n9805, ZN => n9004);
   U2778 : OAI22_X1 port map( A1 => n9262, A2 => n9802, B1 => n2169, B2 => 
                           n9805, ZN => n9005);
   U2779 : OAI22_X1 port map( A1 => n9259, A2 => n9801, B1 => n2161, B2 => 
                           n9804, ZN => n9006);
   U2780 : OAI22_X1 port map( A1 => n9256, A2 => n9802, B1 => n2153, B2 => 
                           n9804, ZN => n9007);
   U2781 : OAI22_X1 port map( A1 => n9253, A2 => n9801, B1 => n2145, B2 => 
                           n9804, ZN => n9008);
   U2782 : OAI22_X1 port map( A1 => n9250, A2 => n9802, B1 => n2137, B2 => 
                           n9804, ZN => n9009);
   U2783 : OAI22_X1 port map( A1 => n9247, A2 => n9801, B1 => n2129, B2 => 
                           n9803, ZN => n9010);
   U2784 : OAI22_X1 port map( A1 => n9244, A2 => n9802, B1 => n2121, B2 => 
                           n9803, ZN => n9011);
   U2785 : OAI22_X1 port map( A1 => n9241, A2 => n9801, B1 => n2113, B2 => 
                           n9803, ZN => n9012);
   U2786 : OAI22_X1 port map( A1 => n9238, A2 => n9802, B1 => n2105, B2 => 
                           n9803, ZN => n9013);
   U2787 : OAI22_X1 port map( A1 => n9331, A2 => n9790, B1 => n2352, B2 => 
                           n9799, ZN => n8950);
   U2788 : OAI22_X1 port map( A1 => n9328, A2 => n9790, B1 => n2344, B2 => 
                           n9799, ZN => n8951);
   U2789 : OAI22_X1 port map( A1 => n9325, A2 => n9790, B1 => n2336, B2 => 
                           n9799, ZN => n8952);
   U2790 : OAI22_X1 port map( A1 => n9322, A2 => n9790, B1 => n2328, B2 => 
                           n9799, ZN => n8953);
   U2791 : OAI22_X1 port map( A1 => n9319, A2 => n9790, B1 => n2320, B2 => 
                           n9798, ZN => n8954);
   U2792 : OAI22_X1 port map( A1 => n9316, A2 => n9790, B1 => n2312, B2 => 
                           n9798, ZN => n8955);
   U2793 : OAI22_X1 port map( A1 => n9313, A2 => n9790, B1 => n2304, B2 => 
                           n9798, ZN => n8956);
   U2794 : OAI22_X1 port map( A1 => n9310, A2 => n9790, B1 => n2296, B2 => 
                           n9798, ZN => n8957);
   U2795 : OAI22_X1 port map( A1 => n9307, A2 => n9790, B1 => n2288, B2 => 
                           n9797, ZN => n8958);
   U2796 : OAI22_X1 port map( A1 => n9304, A2 => n9790, B1 => n2280, B2 => 
                           n9797, ZN => n8959);
   U2797 : OAI22_X1 port map( A1 => n9301, A2 => n9790, B1 => n2272, B2 => 
                           n9797, ZN => n8960);
   U2798 : OAI22_X1 port map( A1 => n9298, A2 => n9790, B1 => n2264, B2 => 
                           n9797, ZN => n8961);
   U2799 : OAI22_X1 port map( A1 => n9295, A2 => n9791, B1 => n2256, B2 => 
                           n9796, ZN => n8962);
   U2800 : OAI22_X1 port map( A1 => n9292, A2 => n9791, B1 => n2248, B2 => 
                           n9796, ZN => n8963);
   U2801 : OAI22_X1 port map( A1 => n9289, A2 => n9791, B1 => n2240, B2 => 
                           n9796, ZN => n8964);
   U2802 : OAI22_X1 port map( A1 => n9286, A2 => n9791, B1 => n2232, B2 => 
                           n9796, ZN => n8965);
   U2803 : OAI22_X1 port map( A1 => n9283, A2 => n9791, B1 => n2224, B2 => 
                           n9795, ZN => n8966);
   U2804 : OAI22_X1 port map( A1 => n9280, A2 => n9791, B1 => n2216, B2 => 
                           n9795, ZN => n8967);
   U2805 : OAI22_X1 port map( A1 => n9277, A2 => n9791, B1 => n2208, B2 => 
                           n9795, ZN => n8968);
   U2806 : OAI22_X1 port map( A1 => n9274, A2 => n9791, B1 => n2200, B2 => 
                           n9795, ZN => n8969);
   U2807 : OAI22_X1 port map( A1 => n9271, A2 => n9791, B1 => n2192, B2 => 
                           n9794, ZN => n8970);
   U2808 : OAI22_X1 port map( A1 => n9268, A2 => n9791, B1 => n2184, B2 => 
                           n9794, ZN => n8971);
   U2809 : OAI22_X1 port map( A1 => n9265, A2 => n9791, B1 => n2176, B2 => 
                           n9794, ZN => n8972);
   U2810 : OAI22_X1 port map( A1 => n9262, A2 => n9791, B1 => n2168, B2 => 
                           n9794, ZN => n8973);
   U2811 : OAI22_X1 port map( A1 => n9259, A2 => n9790, B1 => n2160, B2 => 
                           n9793, ZN => n8974);
   U2812 : OAI22_X1 port map( A1 => n9256, A2 => n9791, B1 => n2152, B2 => 
                           n9793, ZN => n8975);
   U2813 : OAI22_X1 port map( A1 => n9253, A2 => n9790, B1 => n2144, B2 => 
                           n9793, ZN => n8976);
   U2814 : OAI22_X1 port map( A1 => n9250, A2 => n9791, B1 => n2136, B2 => 
                           n9793, ZN => n8977);
   U2815 : OAI22_X1 port map( A1 => n9247, A2 => n9790, B1 => n2128, B2 => 
                           n9792, ZN => n8978);
   U2816 : OAI22_X1 port map( A1 => n9244, A2 => n9791, B1 => n2120, B2 => 
                           n9792, ZN => n8979);
   U2817 : OAI22_X1 port map( A1 => n9241, A2 => n9790, B1 => n2112, B2 => 
                           n9792, ZN => n8980);
   U2818 : OAI22_X1 port map( A1 => n9238, A2 => n9791, B1 => n2104, B2 => 
                           n9792, ZN => n8981);
   U2819 : NAND2_X1 port map( A1 => n1638, A2 => n1639, ZN => OUT2(24));
   U2820 : NOR4_X1 port map( A1 => n1648, A2 => n1649, A3 => n1650, A4 => n1651
                           , ZN => n1638);
   U2821 : NAND2_X1 port map( A1 => n1620, A2 => n1621, ZN => OUT2(25));
   U2822 : NOR4_X1 port map( A1 => n1630, A2 => n1631, A3 => n1632, A4 => n1633
                           , ZN => n1620);
   U2823 : NAND2_X1 port map( A1 => n1602, A2 => n1603, ZN => OUT2(26));
   U2824 : NOR4_X1 port map( A1 => n1612, A2 => n1613, A3 => n1614, A4 => n1615
                           , ZN => n1602);
   U2825 : NAND2_X1 port map( A1 => n1584, A2 => n1585, ZN => OUT2(27));
   U2826 : NOR4_X1 port map( A1 => n1594, A2 => n1595, A3 => n1596, A4 => n1597
                           , ZN => n1584);
   U2827 : NAND2_X1 port map( A1 => n1566, A2 => n1567, ZN => OUT2(28));
   U2828 : NOR4_X1 port map( A1 => n1576, A2 => n1577, A3 => n1578, A4 => n1579
                           , ZN => n1566);
   U2829 : NAND2_X1 port map( A1 => n1548, A2 => n1549, ZN => OUT2(29));
   U2830 : NOR4_X1 port map( A1 => n1558, A2 => n1559, A3 => n1560, A4 => n1561
                           , ZN => n1548);
   U2831 : NAND2_X1 port map( A1 => n1530, A2 => n1531, ZN => OUT2(30));
   U2832 : NOR4_X1 port map( A1 => n1540, A2 => n1541, A3 => n1542, A4 => n1543
                           , ZN => n1530);
   U2833 : NAND2_X1 port map( A1 => n1480, A2 => n1481, ZN => OUT2(31));
   U2834 : NOR4_X1 port map( A1 => n1506, A2 => n1507, A3 => n1508, A4 => n1509
                           , ZN => n1480);
   U2835 : NOR4_X1 port map( A1 => n862, A2 => n863, A3 => n864, A4 => n865, ZN
                           => n861);
   U2836 : OAI221_X1 port map( B1 => n2103, B2 => n9489, C1 => n8406, C2 => 
                           n9486, A => n883, ZN => n862);
   U2837 : NOR4_X1 port map( A1 => n948, A2 => n949, A3 => n950, A4 => n951, ZN
                           => n947);
   U2838 : OAI221_X1 port map( B1 => n2127, B2 => n9489, C1 => n8403, C2 => 
                           n9486, A => n955, ZN => n948);
   U2839 : NOR4_X1 port map( A1 => n1020, A2 => n1021, A3 => n1022, A4 => n1023
                           , ZN => n1019);
   U2840 : OAI221_X1 port map( B1 => n2159, B2 => n9489, C1 => n8399, C2 => 
                           n9486, A => n1027, ZN => n1020);
   U2841 : NOR4_X1 port map( A1 => n1398, A2 => n1399, A3 => n1400, A4 => n1401
                           , ZN => n1397);
   U2842 : OAI221_X1 port map( B1 => n8474, B2 => n9511, C1 => n8238, C2 => 
                           n9508, A => n1403, ZN => n1400);
   U2843 : NOR4_X1 port map( A1 => n1200, A2 => n1201, A3 => n1202, A4 => n1203
                           , ZN => n1199);
   U2844 : OAI221_X1 port map( B1 => n8253, B2 => n9512, C1 => n8216, C2 => 
                           n9509, A => n1205, ZN => n1202);
   U2845 : NOR4_X1 port map( A1 => n1272, A2 => n1273, A3 => n1274, A4 => n1275
                           , ZN => n1271);
   U2846 : OAI221_X1 port map( B1 => n8249, B2 => n9511, C1 => n8224, C2 => 
                           n9508, A => n1277, ZN => n1274);
   U2847 : NOR4_X1 port map( A1 => n1128, A2 => n1129, A3 => n1130, A4 => n1131
                           , ZN => n1127);
   U2848 : OAI221_X1 port map( B1 => n8257, B2 => n9512, C1 => n8208, C2 => 
                           n9509, A => n1133, ZN => n1130);
   U2849 : NOR4_X1 port map( A1 => n930, A2 => n931, A3 => n932, A4 => n933, ZN
                           => n929);
   U2850 : OAI221_X1 port map( B1 => n2119, B2 => n9489, C1 => n8404, C2 => 
                           n9486, A => n937, ZN => n930);
   U2851 : AND3_X1 port map( A1 => ADD_RD2(1), A2 => n10664, A3 => ADD_RD2(2), 
                           ZN => n2079);
   U2852 : AND3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(0), A3 => 
                           ADD_RD2(2), ZN => n2078);
   U2853 : INV_X1 port map( A => ADD_WR(0), ZN => n9921);
   U2854 : INV_X1 port map( A => ADD_WR(2), ZN => n9919);
   U2855 : INV_X1 port map( A => ADD_WR(1), ZN => n9920);
   U2856 : NOR4_X1 port map( A1 => n1344, A2 => n1345, A3 => n1346, A4 => n1347
                           , ZN => n1343);
   U2857 : OAI221_X1 port map( B1 => n8924, B2 => n9439, C1 => n8892, C2 => 
                           n9436, A => n1359, ZN => n1352);
   U2858 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => n10659, A3 => ADD_RD1(2), 
                           ZN => n1467);
   U2859 : INV_X1 port map( A => ADD_RD2(1), ZN => n10663);
   U2860 : INV_X1 port map( A => ADD_RD2(0), ZN => n10664);
   U2861 : NOR4_X1 port map( A1 => n1074, A2 => n1075, A3 => n1076, A4 => n1077
                           , ZN => n1073);
   U2862 : NOR4_X1 port map( A1 => n1082, A2 => n1083, A3 => n1084, A4 => n1085
                           , ZN => n1072);
   U2863 : OAI221_X1 port map( B1 => n8260, B2 => n9512, C1 => n8202, C2 => 
                           n9509, A => n1079, ZN => n1076);
   U2864 : NOR4_X1 port map( A1 => n1326, A2 => n1327, A3 => n1328, A4 => n1329
                           , ZN => n1325);
   U2865 : NOR4_X1 port map( A1 => n1334, A2 => n1335, A3 => n1336, A4 => n1337
                           , ZN => n1324);
   U2866 : OAI221_X1 port map( B1 => n8246, B2 => n9511, C1 => n8230, C2 => 
                           n9508, A => n1331, ZN => n1328);
   U2867 : NOR4_X1 port map( A1 => n1092, A2 => n1093, A3 => n1094, A4 => n1095
                           , ZN => n1091);
   U2868 : NOR4_X1 port map( A1 => n1100, A2 => n1101, A3 => n1102, A4 => n1103
                           , ZN => n1090);
   U2869 : OAI221_X1 port map( B1 => n8259, B2 => n9512, C1 => n8204, C2 => 
                           n9509, A => n1097, ZN => n1094);
   U2870 : AND3_X1 port map( A1 => n10664, A2 => n10663, A3 => ADD_RD2(2), ZN 
                           => n2081);
   U2871 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => n10663, A3 => ADD_RD2(2), 
                           ZN => n2080);
   U2872 : AND3_X1 port map( A1 => n10660, A2 => n10659, A3 => ADD_RD1(2), ZN 
                           => n1466);
   U2873 : NAND2_X1 port map( A1 => n1000, A2 => n1001, ZN => OUT1(25));
   U2874 : NOR4_X1 port map( A1 => n1002, A2 => n1003, A3 => n1004, A4 => n1005
                           , ZN => n1001);
   U2875 : NOR4_X1 port map( A1 => n1010, A2 => n1011, A3 => n1012, A4 => n1013
                           , ZN => n1000);
   U2876 : OAI221_X1 port map( B1 => n2151, B2 => n9489, C1 => n8400, C2 => 
                           n9486, A => n1009, ZN => n1002);
   U2877 : NAND2_X1 port map( A1 => n1378, A2 => n1379, ZN => OUT1(4));
   U2878 : NOR4_X1 port map( A1 => n1380, A2 => n1381, A3 => n1382, A4 => n1383
                           , ZN => n1379);
   U2879 : NOR4_X1 port map( A1 => n1388, A2 => n1389, A3 => n1390, A4 => n1391
                           , ZN => n1378);
   U2880 : OAI221_X1 port map( B1 => n8475, B2 => n9511, C1 => n8236, C2 => 
                           n9508, A => n1385, ZN => n1382);
   U2881 : NAND2_X1 port map( A1 => n1180, A2 => n1181, ZN => OUT1(15));
   U2882 : NOR4_X1 port map( A1 => n1182, A2 => n1183, A3 => n1184, A4 => n1185
                           , ZN => n1181);
   U2883 : NOR4_X1 port map( A1 => n1190, A2 => n1191, A3 => n1192, A4 => n1193
                           , ZN => n1180);
   U2884 : OAI221_X1 port map( B1 => n8254, B2 => n9512, C1 => n8214, C2 => 
                           n9509, A => n1187, ZN => n1184);
   U2885 : NAND2_X1 port map( A1 => n1252, A2 => n1253, ZN => OUT1(11));
   U2886 : NOR4_X1 port map( A1 => n1254, A2 => n1255, A3 => n1256, A4 => n1257
                           , ZN => n1253);
   U2887 : NOR4_X1 port map( A1 => n1262, A2 => n1263, A3 => n1264, A4 => n1265
                           , ZN => n1252);
   U2888 : OAI221_X1 port map( B1 => n8250, B2 => n9511, C1 => n8222, C2 => 
                           n9508, A => n1259, ZN => n1256);
   U2889 : NAND2_X1 port map( A1 => n1108, A2 => n1109, ZN => OUT1(19));
   U2890 : NOR4_X1 port map( A1 => n1110, A2 => n1111, A3 => n1112, A4 => n1113
                           , ZN => n1109);
   U2891 : NOR4_X1 port map( A1 => n1118, A2 => n1119, A3 => n1120, A4 => n1121
                           , ZN => n1108);
   U2892 : OAI221_X1 port map( B1 => n8258, B2 => n9512, C1 => n8206, C2 => 
                           n9509, A => n1115, ZN => n1112);
   U2893 : NAND2_X1 port map( A1 => n1414, A2 => n1415, ZN => OUT1(2));
   U2894 : NOR4_X1 port map( A1 => n1416, A2 => n1417, A3 => n1418, A4 => n1419
                           , ZN => n1415);
   U2895 : NOR4_X1 port map( A1 => n1424, A2 => n1425, A3 => n1426, A4 => n1427
                           , ZN => n1414);
   U2896 : OAI221_X1 port map( B1 => n8473, B2 => n9511, C1 => n8240, C2 => 
                           n9508, A => n1421, ZN => n1418);
   U2897 : NAND2_X1 port map( A1 => n1360, A2 => n1361, ZN => OUT1(5));
   U2898 : NOR4_X1 port map( A1 => n1362, A2 => n1363, A3 => n1364, A4 => n1365
                           , ZN => n1361);
   U2899 : NOR4_X1 port map( A1 => n1370, A2 => n1371, A3 => n1372, A4 => n1373
                           , ZN => n1360);
   U2900 : OAI221_X1 port map( B1 => n8476, B2 => n9511, C1 => n8234, C2 => 
                           n9508, A => n1367, ZN => n1364);
   U2901 : NAND2_X1 port map( A1 => n1162, A2 => n1163, ZN => OUT1(16));
   U2902 : NOR4_X1 port map( A1 => n1164, A2 => n1165, A3 => n1166, A4 => n1167
                           , ZN => n1163);
   U2903 : NOR4_X1 port map( A1 => n1172, A2 => n1173, A3 => n1174, A4 => n1175
                           , ZN => n1162);
   U2904 : OAI221_X1 port map( B1 => n8255, B2 => n9512, C1 => n8212, C2 => 
                           n9509, A => n1169, ZN => n1166);
   U2905 : NAND2_X1 port map( A1 => n1234, A2 => n1235, ZN => OUT1(12));
   U2906 : NOR4_X1 port map( A1 => n1236, A2 => n1237, A3 => n1238, A4 => n1239
                           , ZN => n1235);
   U2907 : NOR4_X1 port map( A1 => n1244, A2 => n1245, A3 => n1246, A4 => n1247
                           , ZN => n1234);
   U2908 : OAI221_X1 port map( B1 => n8251, B2 => n9512, C1 => n8220, C2 => 
                           n9509, A => n1241, ZN => n1238);
   U2909 : NAND2_X1 port map( A1 => n1432, A2 => n1433, ZN => OUT1(1));
   U2910 : NOR4_X1 port map( A1 => n1434, A2 => n1435, A3 => n1436, A4 => n1437
                           , ZN => n1433);
   U2911 : NOR4_X1 port map( A1 => n1442, A2 => n1443, A3 => n1444, A4 => n1445
                           , ZN => n1432);
   U2912 : OAI221_X1 port map( B1 => n8472, B2 => n9511, C1 => n8242, C2 => 
                           n9508, A => n1439, ZN => n1436);
   U2913 : NAND2_X1 port map( A1 => n910, A2 => n911, ZN => OUT1(30));
   U2914 : NOR4_X1 port map( A1 => n912, A2 => n913, A3 => n914, A4 => n915, ZN
                           => n911);
   U2915 : NOR4_X1 port map( A1 => n920, A2 => n921, A3 => n922, A4 => n923, ZN
                           => n910);
   U2916 : OAI221_X1 port map( B1 => n2111, B2 => n9489, C1 => n8405, C2 => 
                           n9486, A => n919, ZN => n912);
   U2917 : NAND2_X1 port map( A1 => n964, A2 => n965, ZN => OUT1(27));
   U2918 : NOR4_X1 port map( A1 => n966, A2 => n967, A3 => n968, A4 => n969, ZN
                           => n965);
   U2919 : NOR4_X1 port map( A1 => n974, A2 => n975, A3 => n976, A4 => n977, ZN
                           => n964);
   U2920 : OAI221_X1 port map( B1 => n2135, B2 => n9489, C1 => n8402, C2 => 
                           n9486, A => n973, ZN => n966);
   U2921 : NAND2_X1 port map( A1 => n1036, A2 => n1037, ZN => OUT1(23));
   U2922 : NOR4_X1 port map( A1 => n1038, A2 => n1039, A3 => n1040, A4 => n1041
                           , ZN => n1037);
   U2923 : NOR4_X1 port map( A1 => n1046, A2 => n1047, A3 => n1048, A4 => n1049
                           , ZN => n1036);
   U2924 : OAI221_X1 port map( B1 => n8262, B2 => n9512, C1 => n8198, C2 => 
                           n9509, A => n1043, ZN => n1040);
   U2925 : NAND2_X1 port map( A1 => n1288, A2 => n1289, ZN => OUT1(9));
   U2926 : NOR4_X1 port map( A1 => n1290, A2 => n1291, A3 => n1292, A4 => n1293
                           , ZN => n1289);
   U2927 : NOR4_X1 port map( A1 => n1298, A2 => n1299, A3 => n1300, A4 => n1301
                           , ZN => n1288);
   U2928 : OAI221_X1 port map( B1 => n8248, B2 => n9511, C1 => n8226, C2 => 
                           n9508, A => n1295, ZN => n1292);
   U2929 : NAND2_X1 port map( A1 => n1054, A2 => n1055, ZN => OUT1(22));
   U2930 : NOR4_X1 port map( A1 => n1056, A2 => n1057, A3 => n1058, A4 => n1059
                           , ZN => n1055);
   U2931 : NOR4_X1 port map( A1 => n1064, A2 => n1065, A3 => n1066, A4 => n1067
                           , ZN => n1054);
   U2932 : OAI221_X1 port map( B1 => n8261, B2 => n9512, C1 => n8200, C2 => 
                           n9509, A => n1061, ZN => n1058);
   U2933 : AND3_X1 port map( A1 => ENABLE, A2 => n9879, A3 => WR, ZN => n849);
   U2934 : INV_X1 port map( A => ADD_RD1(0), ZN => n10660);
   U2935 : NAND2_X1 port map( A1 => n2070, A2 => n2071, ZN => OUT2(0));
   U2936 : NOR4_X1 port map( A1 => n2072, A2 => n2073, A3 => n2074, A4 => n2075
                           , ZN => n2071);
   U2937 : NAND2_X1 port map( A1 => n2052, A2 => n2053, ZN => OUT2(1));
   U2938 : NOR4_X1 port map( A1 => n2054, A2 => n2055, A3 => n2056, A4 => n2057
                           , ZN => n2053);
   U2939 : NAND2_X1 port map( A1 => n2034, A2 => n2035, ZN => OUT2(2));
   U2940 : NOR4_X1 port map( A1 => n2036, A2 => n2037, A3 => n2038, A4 => n2039
                           , ZN => n2035);
   U2941 : NAND2_X1 port map( A1 => n2016, A2 => n2017, ZN => OUT2(3));
   U2942 : NOR4_X1 port map( A1 => n2018, A2 => n2019, A3 => n2020, A4 => n2021
                           , ZN => n2017);
   U2943 : NAND2_X1 port map( A1 => n1998, A2 => n1999, ZN => OUT2(4));
   U2944 : NOR4_X1 port map( A1 => n2000, A2 => n2001, A3 => n2002, A4 => n2003
                           , ZN => n1999);
   U2945 : NAND2_X1 port map( A1 => n1980, A2 => n1981, ZN => OUT2(5));
   U2946 : NOR4_X1 port map( A1 => n1982, A2 => n1983, A3 => n1984, A4 => n1985
                           , ZN => n1981);
   U2947 : NAND2_X1 port map( A1 => n1962, A2 => n1963, ZN => OUT2(6));
   U2948 : NOR4_X1 port map( A1 => n1964, A2 => n1965, A3 => n1966, A4 => n1967
                           , ZN => n1963);
   U2949 : INV_X1 port map( A => DATAIN(3), ZN => n9913);
   U2950 : INV_X1 port map( A => DATAIN(4), ZN => n9912);
   U2951 : INV_X1 port map( A => DATAIN(5), ZN => n9911);
   U2952 : INV_X1 port map( A => DATAIN(6), ZN => n9910);
   U2953 : INV_X1 port map( A => DATAIN(7), ZN => n9909);
   U2954 : INV_X1 port map( A => DATAIN(8), ZN => n9908);
   U2955 : INV_X1 port map( A => DATAIN(31), ZN => n9885);
   U2956 : INV_X1 port map( A => DATAIN(0), ZN => n9916);
   U2957 : INV_X1 port map( A => DATAIN(1), ZN => n9915);
   U2958 : INV_X1 port map( A => DATAIN(2), ZN => n9914);
   U2959 : INV_X1 port map( A => DATAIN(10), ZN => n9906);
   U2960 : INV_X1 port map( A => DATAIN(11), ZN => n9905);
   U2961 : INV_X1 port map( A => DATAIN(12), ZN => n9904);
   U2962 : INV_X1 port map( A => DATAIN(13), ZN => n9903);
   U2963 : INV_X1 port map( A => DATAIN(14), ZN => n9902);
   U2964 : INV_X1 port map( A => DATAIN(15), ZN => n9901);
   U2965 : INV_X1 port map( A => DATAIN(16), ZN => n9900);
   U2966 : INV_X1 port map( A => DATAIN(17), ZN => n9899);
   U2967 : INV_X1 port map( A => DATAIN(18), ZN => n9898);
   U2968 : INV_X1 port map( A => DATAIN(19), ZN => n9897);
   U2969 : INV_X1 port map( A => DATAIN(20), ZN => n9896);
   U2970 : INV_X1 port map( A => DATAIN(21), ZN => n9895);
   U2971 : INV_X1 port map( A => DATAIN(22), ZN => n9894);
   U2972 : INV_X1 port map( A => DATAIN(23), ZN => n9893);
   U2973 : INV_X1 port map( A => DATAIN(24), ZN => n9892);
   U2974 : INV_X1 port map( A => DATAIN(25), ZN => n9891);
   U2975 : INV_X1 port map( A => DATAIN(26), ZN => n9890);
   U2976 : INV_X1 port map( A => DATAIN(27), ZN => n9889);
   U2977 : INV_X1 port map( A => DATAIN(28), ZN => n9888);
   U2978 : INV_X1 port map( A => DATAIN(29), ZN => n9887);
   U2979 : INV_X1 port map( A => DATAIN(30), ZN => n9886);
   U2980 : INV_X1 port map( A => DATAIN(9), ZN => n9907);
   U2981 : INV_X1 port map( A => ADD_RD2(3), ZN => n10662);
   U2982 : INV_X1 port map( A => ADD_RD2(4), ZN => n10661);
   U2983 : INV_X1 port map( A => ADD_RD1(3), ZN => n10658);
   U2984 : NAND2_X1 port map( A1 => n1944, A2 => n1945, ZN => OUT2(7));
   U2985 : NOR4_X1 port map( A1 => n1946, A2 => n1947, A3 => n1948, A4 => n1949
                           , ZN => n1945);
   U2986 : NAND2_X1 port map( A1 => n1926, A2 => n1927, ZN => OUT2(8));
   U2987 : NOR4_X1 port map( A1 => n1936, A2 => n1937, A3 => n1938, A4 => n1939
                           , ZN => n1926);
   U2988 : NAND2_X1 port map( A1 => n1908, A2 => n1909, ZN => OUT2(9));
   U2989 : NOR4_X1 port map( A1 => n1918, A2 => n1919, A3 => n1920, A4 => n1921
                           , ZN => n1908);
   U2990 : NAND2_X1 port map( A1 => n1890, A2 => n1891, ZN => OUT2(10));
   U2991 : NOR4_X1 port map( A1 => n1900, A2 => n1901, A3 => n1902, A4 => n1903
                           , ZN => n1890);
   U2992 : NAND2_X1 port map( A1 => n1872, A2 => n1873, ZN => OUT2(11));
   U2993 : NOR4_X1 port map( A1 => n1882, A2 => n1883, A3 => n1884, A4 => n1885
                           , ZN => n1872);
   U2994 : NAND2_X1 port map( A1 => n1854, A2 => n1855, ZN => OUT2(12));
   U2995 : NOR4_X1 port map( A1 => n1864, A2 => n1865, A3 => n1866, A4 => n1867
                           , ZN => n1854);
   U2996 : NAND2_X1 port map( A1 => n1836, A2 => n1837, ZN => OUT2(13));
   U2997 : NOR4_X1 port map( A1 => n1846, A2 => n1847, A3 => n1848, A4 => n1849
                           , ZN => n1836);
   U2998 : NAND2_X1 port map( A1 => n1818, A2 => n1819, ZN => OUT2(14));
   U2999 : NOR4_X1 port map( A1 => n1828, A2 => n1829, A3 => n1830, A4 => n1831
                           , ZN => n1818);
   U3000 : NAND2_X1 port map( A1 => n1800, A2 => n1801, ZN => OUT2(15));
   U3001 : NOR4_X1 port map( A1 => n1810, A2 => n1811, A3 => n1812, A4 => n1813
                           , ZN => n1800);
   U3002 : NAND2_X1 port map( A1 => n1782, A2 => n1783, ZN => OUT2(16));
   U3003 : NOR4_X1 port map( A1 => n1792, A2 => n1793, A3 => n1794, A4 => n1795
                           , ZN => n1782);
   U3004 : NAND2_X1 port map( A1 => n1764, A2 => n1765, ZN => OUT2(17));
   U3005 : NOR4_X1 port map( A1 => n1774, A2 => n1775, A3 => n1776, A4 => n1777
                           , ZN => n1764);
   U3006 : NAND2_X1 port map( A1 => n1746, A2 => n1747, ZN => OUT2(18));
   U3007 : NOR4_X1 port map( A1 => n1756, A2 => n1757, A3 => n1758, A4 => n1759
                           , ZN => n1746);
   U3008 : NAND2_X1 port map( A1 => n1728, A2 => n1729, ZN => OUT2(19));
   U3009 : NOR4_X1 port map( A1 => n1738, A2 => n1739, A3 => n1740, A4 => n1741
                           , ZN => n1728);
   U3010 : NAND2_X1 port map( A1 => n1710, A2 => n1711, ZN => OUT2(20));
   U3011 : NOR4_X1 port map( A1 => n1720, A2 => n1721, A3 => n1722, A4 => n1723
                           , ZN => n1710);
   U3012 : NAND2_X1 port map( A1 => n1692, A2 => n1693, ZN => OUT2(21));
   U3013 : NOR4_X1 port map( A1 => n1702, A2 => n1703, A3 => n1704, A4 => n1705
                           , ZN => n1692);
   U3014 : NAND2_X1 port map( A1 => n1674, A2 => n1675, ZN => OUT2(22));
   U3015 : NOR4_X1 port map( A1 => n1684, A2 => n1685, A3 => n1686, A4 => n1687
                           , ZN => n1674);
   U3016 : NAND2_X1 port map( A1 => n1656, A2 => n1657, ZN => OUT2(23));
   U3017 : NOR4_X1 port map( A1 => n1666, A2 => n1667, A3 => n1668, A4 => n1669
                           , ZN => n1656);
   U3018 : INV_X1 port map( A => ADD_WR(4), ZN => n9917);
   U3019 : INV_X1 port map( A => ADD_WR(3), ZN => n9918);
   U3020 : OAI221_X1 port map( B1 => n8667, B2 => n9476, C1 => n8643, C2 => 
                           n9473, A => n1230, ZN => n1229);
   U3021 : OAI221_X1 port map( B1 => n8787, B2 => n9464, C1 => n8219, C2 => 
                           n9461, A => n1231, ZN => n1228);
   U3022 : OAI221_X1 port map( B1 => n8671, B2 => n9476, C1 => n8647, C2 => 
                           n9473, A => n1158, ZN => n1157);
   U3023 : OAI221_X1 port map( B1 => n8791, B2 => n9464, C1 => n8211, C2 => 
                           n9461, A => n1159, ZN => n1156);
   U3024 : OAI221_X1 port map( B1 => n8598, B2 => n9523, C1 => n8566, C2 => 
                           n9520, A => n1456, ZN => n1455);
   U3025 : AOI22_X1 port map( A1 => n9517, A2 => n10473, B1 => n9516, B2 => 
                           n10289, ZN => n1456);
   U3026 : NAND2_X1 port map( A1 => n1270, A2 => n1271, ZN => OUT1(10));
   U3027 : NOR4_X1 port map( A1 => n1280, A2 => n1281, A3 => n1282, A4 => n1283
                           , ZN => n1270);
   U3028 : NAND2_X1 port map( A1 => n928, A2 => n929, ZN => OUT1(29));
   U3029 : NOR4_X1 port map( A1 => n938, A2 => n939, A3 => n940, A4 => n941, ZN
                           => n928);
   U3030 : NAND2_X1 port map( A1 => n1324, A2 => n1325, ZN => OUT1(7));
   U3031 : NAND2_X1 port map( A1 => n1018, A2 => n1019, ZN => OUT1(24));
   U3032 : NOR4_X1 port map( A1 => n1028, A2 => n1029, A3 => n1030, A4 => n1031
                           , ZN => n1018);
   U3033 : NAND2_X1 port map( A1 => n1090, A2 => n1091, ZN => OUT1(20));
   U3034 : NAND2_X1 port map( A1 => n1072, A2 => n1073, ZN => OUT1(21));
   U3035 : OAI221_X1 port map( B1 => n8654, B2 => n9475, C1 => n8630, C2 => 
                           n9472, A => n1475, ZN => n1474);
   U3036 : OAI221_X1 port map( B1 => n8774, B2 => n9463, C1 => n8245, C2 => 
                           n9460, A => n1476, ZN => n1473);
   U3037 : NAND2_X1 port map( A1 => n1198, A2 => n1199, ZN => OUT1(14));
   U3038 : NOR4_X1 port map( A1 => n1208, A2 => n1209, A3 => n1210, A4 => n1211
                           , ZN => n1198);
   U3039 : NAND2_X1 port map( A1 => n1126, A2 => n1127, ZN => OUT1(18));
   U3040 : NOR4_X1 port map( A1 => n1136, A2 => n1137, A3 => n1138, A4 => n1139
                           , ZN => n1126);
   U3041 : NAND2_X1 port map( A1 => n946, A2 => n947, ZN => OUT1(28));
   U3042 : NOR4_X1 port map( A1 => n956, A2 => n957, A3 => n958, A4 => n959, ZN
                           => n946);
   U3043 : NAND2_X1 port map( A1 => n860, A2 => n861, ZN => OUT1(31));
   U3044 : NOR4_X1 port map( A1 => n886, A2 => n887, A3 => n888, A4 => n889, ZN
                           => n860);
   U3045 : NAND2_X1 port map( A1 => n1396, A2 => n1397, ZN => OUT1(3));
   U3046 : NOR4_X1 port map( A1 => n1406, A2 => n1407, A3 => n1408, A4 => n1409
                           , ZN => n1396);
   U3047 : NAND2_X1 port map( A1 => n1216, A2 => n1217, ZN => OUT1(13));
   U3048 : NOR4_X1 port map( A1 => n1226, A2 => n1227, A3 => n1228, A4 => n1229
                           , ZN => n1216);
   U3049 : NAND2_X1 port map( A1 => n1144, A2 => n1145, ZN => OUT1(17));
   U3050 : NOR4_X1 port map( A1 => n1154, A2 => n1155, A3 => n1156, A4 => n1157
                           , ZN => n1144);
   U3051 : NAND2_X1 port map( A1 => n1450, A2 => n1451, ZN => OUT1(0));
   U3052 : NOR4_X1 port map( A1 => n1471, A2 => n1472, A3 => n1473, A4 => n1474
                           , ZN => n1450);
   U3053 : AND3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(0), A3 => 
                           ADD_RD1(2), ZN => n1464);
   U3054 : AND3_X1 port map( A1 => ADD_RD1(1), A2 => n10660, A3 => ADD_RD1(2), 
                           ZN => n1468);
   U3055 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => 
                           ADD_RD1(0), ZN => n1457);
   U3056 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n10660, 
                           ZN => n1459);
   U3057 : INV_X1 port map( A => ADD_RD1(1), ZN => n10659);
   U3058 : INV_X1 port map( A => ADD_RD1(4), ZN => n10665);
   U3059 : NOR4_X1 port map( A1 => n1352, A2 => n1353, A3 => n1354, A4 => n1355
                           , ZN => n1342);
   U3060 : OAI221_X1 port map( B1 => n8660, B2 => n9475, C1 => n8636, C2 => 
                           n9472, A => n1356, ZN => n1355);
   U3061 : OAI221_X1 port map( B1 => n8780, B2 => n9463, C1 => n8233, C2 => 
                           n9460, A => n1357, ZN => n1354);
   U3062 : NAND2_X1 port map( A1 => n1342, A2 => n1343, ZN => OUT1(6));
   U3063 : NAND2_X1 port map( A1 => n1306, A2 => n1307, ZN => OUT1(8));
   U3064 : CLKBUF_X1 port map( A => n9882, Z => n9877);
   U3065 : CLKBUF_X1 port map( A => n9881, Z => n9878);
   U3066 : CLKBUF_X1 port map( A => n9880, Z => n9879);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_9 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_9;

architecture SYN_behavioral of reg_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n34, n35, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n35, Z => n177);
   U4 : BUF_X1 port map( A => n35, Z => n176);
   U5 : BUF_X1 port map( A => n35, Z => n178);
   U6 : BUF_X1 port map( A => n34, Z => n179);
   U7 : BUF_X1 port map( A => n34, Z => n180);
   U8 : BUF_X1 port map( A => n34, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n35);
   U10 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n190, ZN 
                           => n75);
   U11 : INV_X1 port map( A => i(24), ZN => n190);
   U12 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n189, ZN 
                           => n74);
   U13 : INV_X1 port map( A => i(25), ZN => n189);
   U14 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n188, ZN 
                           => n73);
   U15 : INV_X1 port map( A => i(26), ZN => n188);
   U16 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n187, ZN 
                           => n72);
   U17 : INV_X1 port map( A => i(27), ZN => n187);
   U18 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n186, ZN 
                           => n71);
   U19 : INV_X1 port map( A => i(28), ZN => n186);
   U20 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U21 : INV_X1 port map( A => i(29), ZN => n185);
   U22 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U23 : INV_X1 port map( A => i(30), ZN => n184);
   U24 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U25 : INV_X1 port map( A => i(31), ZN => n183);
   U26 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U27 : INV_X1 port map( A => i(0), ZN => n214);
   U28 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U29 : INV_X1 port map( A => i(1), ZN => n213);
   U30 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U31 : INV_X1 port map( A => i(2), ZN => n212);
   U32 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U33 : INV_X1 port map( A => i(3), ZN => n211);
   U34 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U35 : INV_X1 port map( A => i(4), ZN => n210);
   U36 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U37 : INV_X1 port map( A => i(5), ZN => n209);
   U38 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U39 : INV_X1 port map( A => i(6), ZN => n208);
   U40 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U41 : INV_X1 port map( A => i(7), ZN => n207);
   U42 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U43 : INV_X1 port map( A => i(8), ZN => n206);
   U44 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U45 : INV_X1 port map( A => i(9), ZN => n205);
   U46 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U47 : INV_X1 port map( A => i(10), ZN => n204);
   U48 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U49 : INV_X1 port map( A => i(11), ZN => n203);
   U50 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U51 : INV_X1 port map( A => i(12), ZN => n202);
   U52 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U53 : INV_X1 port map( A => i(13), ZN => n201);
   U54 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U55 : INV_X1 port map( A => i(14), ZN => n200);
   U56 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n199, ZN 
                           => n84);
   U57 : INV_X1 port map( A => i(15), ZN => n199);
   U58 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n198, ZN 
                           => n83);
   U59 : INV_X1 port map( A => i(16), ZN => n198);
   U60 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n197, ZN 
                           => n82);
   U61 : INV_X1 port map( A => i(17), ZN => n197);
   U62 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n196, ZN 
                           => n81);
   U63 : INV_X1 port map( A => i(18), ZN => n196);
   U64 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n195, ZN 
                           => n80);
   U65 : INV_X1 port map( A => i(19), ZN => n195);
   U66 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n194, ZN 
                           => n79);
   U67 : INV_X1 port map( A => i(20), ZN => n194);
   U68 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n193, ZN 
                           => n78);
   U69 : INV_X1 port map( A => i(21), ZN => n193);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n192, ZN 
                           => n77);
   U71 : INV_X1 port map( A => i(22), ZN => n192);
   U72 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n191, ZN 
                           => n76);
   U73 : INV_X1 port map( A => i(23), ZN => n191);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n34);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_10 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_10;

architecture SYN_behavioral of reg_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n34, n35, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n35, Z => n177);
   U4 : BUF_X1 port map( A => n35, Z => n176);
   U5 : BUF_X1 port map( A => n35, Z => n178);
   U6 : BUF_X1 port map( A => n34, Z => n179);
   U7 : BUF_X1 port map( A => n34, Z => n180);
   U8 : BUF_X1 port map( A => n34, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n35);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U11 : INV_X1 port map( A => i(6), ZN => n208);
   U12 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U13 : INV_X1 port map( A => i(12), ZN => n202);
   U14 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n198, ZN 
                           => n83);
   U15 : INV_X1 port map( A => i(16), ZN => n198);
   U16 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n194, ZN 
                           => n79);
   U17 : INV_X1 port map( A => i(20), ZN => n194);
   U18 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n187, ZN 
                           => n72);
   U19 : INV_X1 port map( A => i(27), ZN => n187);
   U20 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U21 : INV_X1 port map( A => i(30), ZN => n184);
   U22 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U23 : INV_X1 port map( A => i(0), ZN => n214);
   U24 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U25 : INV_X1 port map( A => i(13), ZN => n201);
   U26 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n197, ZN 
                           => n82);
   U27 : INV_X1 port map( A => i(17), ZN => n197);
   U28 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n190, ZN 
                           => n75);
   U29 : INV_X1 port map( A => i(24), ZN => n190);
   U30 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n186, ZN 
                           => n71);
   U31 : INV_X1 port map( A => i(28), ZN => n186);
   U32 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U33 : INV_X1 port map( A => i(31), ZN => n183);
   U34 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U35 : INV_X1 port map( A => i(3), ZN => n211);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U37 : INV_X1 port map( A => i(10), ZN => n204);
   U38 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U39 : INV_X1 port map( A => i(14), ZN => n200);
   U40 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n196, ZN 
                           => n81);
   U41 : INV_X1 port map( A => i(18), ZN => n196);
   U42 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U43 : INV_X1 port map( A => i(29), ZN => n185);
   U44 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U45 : INV_X1 port map( A => i(8), ZN => n206);
   U46 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U47 : INV_X1 port map( A => i(7), ZN => n207);
   U48 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n193, ZN 
                           => n78);
   U49 : INV_X1 port map( A => i(21), ZN => n193);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n189, ZN 
                           => n74);
   U51 : INV_X1 port map( A => i(25), ZN => n189);
   U52 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U53 : INV_X1 port map( A => i(2), ZN => n212);
   U54 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U55 : INV_X1 port map( A => i(4), ZN => n210);
   U56 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U57 : INV_X1 port map( A => i(11), ZN => n203);
   U58 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n199, ZN 
                           => n84);
   U59 : INV_X1 port map( A => i(15), ZN => n199);
   U60 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n195, ZN 
                           => n80);
   U61 : INV_X1 port map( A => i(19), ZN => n195);
   U62 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n188, ZN 
                           => n73);
   U63 : INV_X1 port map( A => i(26), ZN => n188);
   U64 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U65 : INV_X1 port map( A => i(1), ZN => n213);
   U66 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U67 : INV_X1 port map( A => i(5), ZN => n209);
   U68 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U69 : INV_X1 port map( A => i(9), ZN => n205);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n191, ZN 
                           => n76);
   U71 : INV_X1 port map( A => i(23), ZN => n191);
   U72 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n192, ZN 
                           => n77);
   U73 : INV_X1 port map( A => i(22), ZN => n192);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n34);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_11 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_11;

architecture SYN_behavioral of reg_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n34, n35, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n35, Z => n177);
   U4 : BUF_X1 port map( A => n35, Z => n176);
   U5 : BUF_X1 port map( A => n35, Z => n178);
   U6 : BUF_X1 port map( A => n34, Z => n179);
   U7 : BUF_X1 port map( A => n34, Z => n180);
   U8 : BUF_X1 port map( A => n34, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n35);
   U10 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U11 : INV_X1 port map( A => i(10), ZN => n204);
   U12 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U13 : INV_X1 port map( A => i(11), ZN => n203);
   U14 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U15 : INV_X1 port map( A => i(12), ZN => n202);
   U16 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U17 : INV_X1 port map( A => i(13), ZN => n201);
   U18 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U19 : INV_X1 port map( A => i(14), ZN => n200);
   U20 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U21 : INV_X1 port map( A => i(0), ZN => n214);
   U22 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U23 : INV_X1 port map( A => i(8), ZN => n206);
   U24 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U25 : INV_X1 port map( A => i(3), ZN => n211);
   U26 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U27 : INV_X1 port map( A => i(4), ZN => n210);
   U28 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U29 : INV_X1 port map( A => i(9), ZN => n205);
   U30 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U31 : INV_X1 port map( A => i(2), ZN => n212);
   U32 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U33 : INV_X1 port map( A => i(5), ZN => n209);
   U34 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U35 : INV_X1 port map( A => i(6), ZN => n208);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U37 : INV_X1 port map( A => i(7), ZN => n207);
   U38 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n185, ZN 
                           => n77);
   U39 : INV_X1 port map( A => i(22), ZN => n185);
   U40 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n193, ZN 
                           => n74);
   U41 : INV_X1 port map( A => i(25), ZN => n193);
   U42 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n194, ZN 
                           => n73);
   U43 : INV_X1 port map( A => i(26), ZN => n194);
   U44 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n195, ZN 
                           => n72);
   U45 : INV_X1 port map( A => i(27), ZN => n195);
   U46 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n196, ZN 
                           => n71);
   U47 : INV_X1 port map( A => i(28), ZN => n196);
   U48 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n197, ZN 
                           => n70);
   U49 : INV_X1 port map( A => i(29), ZN => n197);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n198, ZN 
                           => n69);
   U51 : INV_X1 port map( A => i(30), ZN => n198);
   U52 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n199, ZN 
                           => n68);
   U53 : INV_X1 port map( A => i(31), ZN => n199);
   U54 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n192, ZN 
                           => n84);
   U55 : INV_X1 port map( A => i(15), ZN => n192);
   U56 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n191, ZN 
                           => n83);
   U57 : INV_X1 port map( A => i(16), ZN => n191);
   U58 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n190, ZN 
                           => n82);
   U59 : INV_X1 port map( A => i(17), ZN => n190);
   U60 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n189, ZN 
                           => n81);
   U61 : INV_X1 port map( A => i(18), ZN => n189);
   U62 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n188, ZN 
                           => n80);
   U63 : INV_X1 port map( A => i(19), ZN => n188);
   U64 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n187, ZN 
                           => n79);
   U65 : INV_X1 port map( A => i(20), ZN => n187);
   U66 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n186, ZN 
                           => n78);
   U67 : INV_X1 port map( A => i(21), ZN => n186);
   U68 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n184, ZN 
                           => n76);
   U69 : INV_X1 port map( A => i(23), ZN => n184);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n183, ZN 
                           => n75);
   U71 : INV_X1 port map( A => i(24), ZN => n183);
   U72 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U73 : INV_X1 port map( A => i(1), ZN => n213);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n34);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity BranchUnit is

   port( a : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : out 
         std_logic);

end BranchUnit;

architecture SYN_Behavioral of BranchUnit is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   U2 : NOR4_X1 port map( A1 => a(5), A2 => a(4), A3 => a(3), A4 => a(31), ZN 
                           => n10);
   U3 : NOR4_X1 port map( A1 => a(1), A2 => a(19), A3 => a(18), A4 => a(17), ZN
                           => n6);
   U4 : NOR4_X1 port map( A1 => a(12), A2 => a(11), A3 => a(10), A4 => a(0), ZN
                           => n4);
   U5 : NOR4_X1 port map( A1 => a(16), A2 => a(15), A3 => a(14), A4 => a(13), 
                           ZN => n5);
   U6 : NOR4_X1 port map( A1 => a(30), A2 => a(2), A3 => a(29), A4 => a(28), ZN
                           => n9);
   U7 : NOR4_X1 port map( A1 => a(27), A2 => a(26), A3 => a(25), A4 => a(24), 
                           ZN => n8);
   U8 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => n1);
   U9 : NAND4_X1 port map( A1 => n8, A2 => n9, A3 => n10, A4 => n11, ZN => n2);
   U10 : NOR4_X1 port map( A1 => a(9), A2 => a(8), A3 => a(7), A4 => a(6), ZN 
                           => n11);
   U11 : NAND4_X1 port map( A1 => n4, A2 => n5, A3 => n6, A4 => n7, ZN => n3);
   U12 : NOR4_X1 port map( A1 => a(23), A2 => a(22), A3 => a(21), A4 => a(20), 
                           ZN => n7);
   U13 : XNOR2_X1 port map( A => sel, B => n1, ZN => y);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Mux21_5 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end Mux21_5;

architecture SYN_Behavioral of Mux21_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n148, Z => n140);
   U2 : BUF_X1 port map( A => n145, Z => n147);
   U3 : BUF_X1 port map( A => n143, Z => n146);
   U4 : BUF_X1 port map( A => n148, Z => n145);
   U5 : BUF_X1 port map( A => n148, Z => n144);
   U6 : BUF_X1 port map( A => n148, Z => n141);
   U7 : BUF_X1 port map( A => n148, Z => n143);
   U8 : BUF_X1 port map( A => n148, Z => n142);
   U9 : INV_X1 port map( A => n139, ZN => n148);
   U10 : INV_X1 port map( A => n38, ZN => y(5));
   U11 : AOI22_X1 port map( A1 => a(5), A2 => sel, B1 => b(5), B2 => n141, ZN 
                           => n38);
   U12 : INV_X1 port map( A => n37, ZN => y(6));
   U13 : AOI22_X1 port map( A1 => a(6), A2 => n139, B1 => b(6), B2 => n140, ZN 
                           => n37);
   U14 : INV_X1 port map( A => n62, ZN => y(12));
   U15 : AOI22_X1 port map( A1 => a(12), A2 => sel, B1 => b(12), B2 => n147, ZN
                           => n62);
   U16 : INV_X1 port map( A => n61, ZN => y(13));
   U17 : AOI22_X1 port map( A1 => a(13), A2 => n139, B1 => b(13), B2 => n146, 
                           ZN => n61);
   U18 : INV_X1 port map( A => n60, ZN => y(14));
   U19 : AOI22_X1 port map( A1 => a(14), A2 => sel, B1 => b(14), B2 => n146, ZN
                           => n60);
   U20 : INV_X1 port map( A => n34, ZN => y(9));
   U21 : AOI22_X1 port map( A1 => n139, A2 => a(9), B1 => b(9), B2 => n140, ZN 
                           => n34);
   U22 : INV_X1 port map( A => n35, ZN => y(8));
   U23 : AOI22_X1 port map( A1 => a(8), A2 => sel, B1 => b(8), B2 => n140, ZN 
                           => n35);
   U24 : INV_X1 port map( A => n39, ZN => y(4));
   U25 : AOI22_X1 port map( A1 => a(4), A2 => n139, B1 => b(4), B2 => n141, ZN 
                           => n39);
   U26 : INV_X1 port map( A => n40, ZN => y(3));
   U27 : AOI22_X1 port map( A1 => a(3), A2 => sel, B1 => b(3), B2 => n141, ZN 
                           => n40);
   U28 : INV_X1 port map( A => n43, ZN => y(2));
   U29 : AOI22_X1 port map( A1 => a(2), A2 => sel, B1 => b(2), B2 => n142, ZN 
                           => n43);
   U30 : INV_X1 port map( A => n36, ZN => y(7));
   U31 : AOI22_X1 port map( A1 => a(7), A2 => n139, B1 => b(7), B2 => n140, ZN 
                           => n36);
   U32 : INV_X1 port map( A => n64, ZN => y(10));
   U33 : AOI22_X1 port map( A1 => a(10), A2 => n139, B1 => b(10), B2 => n147, 
                           ZN => n64);
   U34 : INV_X1 port map( A => n63, ZN => y(11));
   U35 : AOI22_X1 port map( A1 => a(11), A2 => sel, B1 => b(11), B2 => n147, ZN
                           => n63);
   U36 : INV_X1 port map( A => n65, ZN => y(0));
   U37 : AOI22_X1 port map( A1 => a(0), A2 => n139, B1 => b(0), B2 => n147, ZN 
                           => n65);
   U38 : INV_X1 port map( A => n51, ZN => y(22));
   U39 : INV_X1 port map( A => n48, ZN => y(25));
   U40 : INV_X1 port map( A => n47, ZN => y(26));
   U41 : INV_X1 port map( A => n46, ZN => y(27));
   U42 : INV_X1 port map( A => n45, ZN => y(28));
   U43 : INV_X1 port map( A => n44, ZN => y(29));
   U44 : INV_X1 port map( A => n42, ZN => y(30));
   U45 : INV_X1 port map( A => n41, ZN => y(31));
   U46 : INV_X1 port map( A => n59, ZN => y(15));
   U47 : AOI22_X1 port map( A1 => a(15), A2 => sel, B1 => b(15), B2 => n146, ZN
                           => n59);
   U48 : INV_X1 port map( A => n58, ZN => y(16));
   U49 : AOI22_X1 port map( A1 => a(16), A2 => n139, B1 => b(16), B2 => n146, 
                           ZN => n58);
   U50 : INV_X1 port map( A => n57, ZN => y(17));
   U51 : AOI22_X1 port map( A1 => a(17), A2 => sel, B1 => b(17), B2 => n145, ZN
                           => n57);
   U52 : INV_X1 port map( A => n56, ZN => y(18));
   U53 : AOI22_X1 port map( A1 => a(18), A2 => n139, B1 => b(18), B2 => n145, 
                           ZN => n56);
   U54 : INV_X1 port map( A => n55, ZN => y(19));
   U55 : AOI22_X1 port map( A1 => a(19), A2 => sel, B1 => b(19), B2 => n145, ZN
                           => n55);
   U56 : INV_X1 port map( A => n53, ZN => y(20));
   U57 : AOI22_X1 port map( A1 => a(20), A2 => n139, B1 => b(20), B2 => n144, 
                           ZN => n53);
   U58 : INV_X1 port map( A => n52, ZN => y(21));
   U59 : AOI22_X1 port map( A1 => a(21), A2 => sel, B1 => b(21), B2 => n144, ZN
                           => n52);
   U60 : INV_X1 port map( A => n50, ZN => y(23));
   U61 : AOI22_X1 port map( A1 => a(23), A2 => n139, B1 => b(23), B2 => n144, 
                           ZN => n50);
   U62 : INV_X1 port map( A => n49, ZN => y(24));
   U63 : AOI22_X1 port map( A1 => a(24), A2 => sel, B1 => b(24), B2 => n143, ZN
                           => n49);
   U64 : INV_X1 port map( A => n54, ZN => y(1));
   U65 : AOI22_X1 port map( A1 => a(1), A2 => n139, B1 => b(1), B2 => n145, ZN 
                           => n54);
   U66 : BUF_X1 port map( A => sel, Z => n139);
   U67 : AOI22_X1 port map( A1 => a(22), A2 => n139, B1 => b(22), B2 => n144, 
                           ZN => n51);
   U68 : AOI22_X1 port map( A1 => a(31), A2 => sel, B1 => b(31), B2 => n141, ZN
                           => n41);
   U69 : AOI22_X1 port map( A1 => a(30), A2 => n139, B1 => b(30), B2 => n142, 
                           ZN => n42);
   U70 : AOI22_X1 port map( A1 => a(29), A2 => sel, B1 => b(29), B2 => n142, ZN
                           => n44);
   U71 : AOI22_X1 port map( A1 => a(28), A2 => n139, B1 => b(28), B2 => n142, 
                           ZN => n45);
   U72 : AOI22_X1 port map( A1 => a(27), A2 => sel, B1 => b(27), B2 => n143, ZN
                           => n46);
   U73 : AOI22_X1 port map( A1 => a(26), A2 => n139, B1 => b(26), B2 => n143, 
                           ZN => n47);
   U74 : AOI22_X1 port map( A1 => a(25), A2 => sel, B1 => b(25), B2 => n143, ZN
                           => n48);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Mux41 is

   port( a, b, c, d : in std_logic_vector (31 downto 0);  sel : in 
         std_logic_vector (1 downto 0);  y : out std_logic_vector (31 downto 0)
         );

end Mux41;

architecture SYN_Behavioral of Mux41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n6, Z => n157);
   U2 : BUF_X1 port map( A => n6, Z => n158);
   U3 : BUF_X1 port map( A => n4, Z => n163);
   U4 : BUF_X1 port map( A => n4, Z => n164);
   U5 : BUF_X1 port map( A => n7, Z => n154);
   U6 : BUF_X1 port map( A => n7, Z => n155);
   U7 : BUF_X1 port map( A => n5, Z => n160);
   U8 : BUF_X1 port map( A => n5, Z => n161);
   U9 : BUF_X1 port map( A => n6, Z => n159);
   U10 : BUF_X1 port map( A => n4, Z => n165);
   U11 : BUF_X1 port map( A => n7, Z => n156);
   U12 : BUF_X1 port map( A => n5, Z => n162);
   U13 : AOI22_X1 port map( A1 => a(4), A2 => n159, B1 => b(4), B2 => n156, ZN 
                           => n16);
   U14 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => y(0));
   U15 : AOI22_X1 port map( A1 => c(0), A2 => n163, B1 => d(0), B2 => n160, ZN 
                           => n69);
   U16 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => y(4));
   U17 : AOI22_X1 port map( A1 => c(4), A2 => n165, B1 => d(4), B2 => n162, ZN 
                           => n17);
   U18 : AOI22_X1 port map( A1 => a(3), A2 => n159, B1 => b(3), B2 => n156, ZN 
                           => n18);
   U19 : AOI22_X1 port map( A1 => a(0), A2 => n157, B1 => b(0), B2 => n154, ZN 
                           => n68);
   U20 : AOI22_X1 port map( A1 => a(1), A2 => n157, B1 => b(1), B2 => n154, ZN 
                           => n46);
   U21 : AOI22_X1 port map( A1 => a(2), A2 => n158, B1 => b(2), B2 => n155, ZN 
                           => n24);
   U22 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => y(2));
   U23 : AOI22_X1 port map( A1 => c(2), A2 => n164, B1 => d(2), B2 => n161, ZN 
                           => n25);
   U24 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => y(1));
   U25 : AOI22_X1 port map( A1 => c(1), A2 => n163, B1 => d(1), B2 => n160, ZN 
                           => n47);
   U26 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => y(3));
   U27 : AOI22_X1 port map( A1 => c(3), A2 => n165, B1 => d(3), B2 => n162, ZN 
                           => n19);
   U28 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => y(5));
   U29 : AOI22_X1 port map( A1 => a(5), A2 => n159, B1 => b(5), B2 => n156, ZN 
                           => n14);
   U30 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => y(6));
   U31 : AOI22_X1 port map( A1 => a(6), A2 => n159, B1 => b(6), B2 => n156, ZN 
                           => n12);
   U32 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => y(20));
   U33 : AOI22_X1 port map( A1 => a(20), A2 => n158, B1 => b(20), B2 => n155, 
                           ZN => n44);
   U34 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => y(21));
   U35 : AOI22_X1 port map( A1 => a(21), A2 => n158, B1 => b(21), B2 => n155, 
                           ZN => n42);
   U36 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => y(22));
   U37 : AOI22_X1 port map( A1 => a(22), A2 => n158, B1 => b(22), B2 => n155, 
                           ZN => n40);
   U38 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => y(23));
   U39 : AOI22_X1 port map( A1 => a(23), A2 => n158, B1 => b(23), B2 => n155, 
                           ZN => n38);
   U40 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => y(24));
   U41 : AOI22_X1 port map( A1 => a(24), A2 => n158, B1 => b(24), B2 => n155, 
                           ZN => n36);
   U42 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => y(25));
   U43 : AOI22_X1 port map( A1 => a(25), A2 => n158, B1 => b(25), B2 => n155, 
                           ZN => n34);
   U44 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => y(26));
   U45 : AOI22_X1 port map( A1 => a(26), A2 => n158, B1 => b(26), B2 => n155, 
                           ZN => n32);
   U46 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => y(27));
   U47 : AOI22_X1 port map( A1 => a(27), A2 => n158, B1 => b(27), B2 => n155, 
                           ZN => n30);
   U48 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => y(28));
   U49 : AOI22_X1 port map( A1 => a(28), A2 => n158, B1 => b(28), B2 => n155, 
                           ZN => n28);
   U50 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => y(29));
   U51 : AOI22_X1 port map( A1 => a(29), A2 => n158, B1 => b(29), B2 => n155, 
                           ZN => n26);
   U52 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => y(30));
   U53 : AOI22_X1 port map( A1 => a(30), A2 => n158, B1 => b(30), B2 => n155, 
                           ZN => n22);
   U54 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => y(31));
   U55 : AOI22_X1 port map( A1 => a(31), A2 => n159, B1 => b(31), B2 => n156, 
                           ZN => n20);
   U56 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => y(7));
   U57 : AOI22_X1 port map( A1 => a(7), A2 => n159, B1 => b(7), B2 => n156, ZN 
                           => n10);
   U58 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => y(8));
   U59 : AOI22_X1 port map( A1 => a(8), A2 => n159, B1 => b(8), B2 => n156, ZN 
                           => n8);
   U60 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => y(9));
   U61 : AOI22_X1 port map( A1 => a(9), A2 => n159, B1 => b(9), B2 => n156, ZN 
                           => n2);
   U62 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => y(10));
   U63 : AOI22_X1 port map( A1 => a(10), A2 => n157, B1 => b(10), B2 => n154, 
                           ZN => n66);
   U64 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => y(11));
   U65 : AOI22_X1 port map( A1 => a(11), A2 => n157, B1 => b(11), B2 => n154, 
                           ZN => n64);
   U66 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => y(12));
   U67 : AOI22_X1 port map( A1 => a(12), A2 => n157, B1 => b(12), B2 => n154, 
                           ZN => n62);
   U68 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => y(13));
   U69 : AOI22_X1 port map( A1 => a(13), A2 => n157, B1 => b(13), B2 => n154, 
                           ZN => n60);
   U70 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => y(14));
   U71 : AOI22_X1 port map( A1 => a(14), A2 => n157, B1 => b(14), B2 => n154, 
                           ZN => n58);
   U72 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => y(15));
   U73 : AOI22_X1 port map( A1 => a(15), A2 => n157, B1 => b(15), B2 => n154, 
                           ZN => n56);
   U74 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => y(16));
   U75 : AOI22_X1 port map( A1 => a(16), A2 => n157, B1 => b(16), B2 => n154, 
                           ZN => n54);
   U76 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => y(17));
   U77 : AOI22_X1 port map( A1 => a(17), A2 => n157, B1 => b(17), B2 => n154, 
                           ZN => n52);
   U78 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => y(18));
   U79 : AOI22_X1 port map( A1 => a(18), A2 => n157, B1 => b(18), B2 => n154, 
                           ZN => n50);
   U80 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => y(19));
   U81 : AOI22_X1 port map( A1 => a(19), A2 => n157, B1 => b(19), B2 => n154, 
                           ZN => n48);
   U82 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n6);
   U83 : NOR2_X1 port map( A1 => n166, A2 => sel(1), ZN => n7);
   U84 : AND2_X1 port map( A1 => sel(1), A2 => n166, ZN => n4);
   U85 : AND2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n5);
   U86 : INV_X1 port map( A => sel(0), ZN => n166);
   U87 : AOI22_X1 port map( A1 => c(5), A2 => n165, B1 => d(5), B2 => n162, ZN 
                           => n15);
   U88 : AOI22_X1 port map( A1 => c(6), A2 => n165, B1 => d(6), B2 => n162, ZN 
                           => n13);
   U89 : AOI22_X1 port map( A1 => c(7), A2 => n165, B1 => d(7), B2 => n162, ZN 
                           => n11);
   U90 : AOI22_X1 port map( A1 => c(8), A2 => n165, B1 => d(8), B2 => n162, ZN 
                           => n9);
   U91 : AOI22_X1 port map( A1 => c(9), A2 => n165, B1 => d(9), B2 => n162, ZN 
                           => n3);
   U92 : AOI22_X1 port map( A1 => c(10), A2 => n163, B1 => d(10), B2 => n160, 
                           ZN => n67);
   U93 : AOI22_X1 port map( A1 => c(11), A2 => n163, B1 => d(11), B2 => n160, 
                           ZN => n65);
   U94 : AOI22_X1 port map( A1 => c(12), A2 => n163, B1 => d(12), B2 => n160, 
                           ZN => n63);
   U95 : AOI22_X1 port map( A1 => c(13), A2 => n163, B1 => d(13), B2 => n160, 
                           ZN => n61);
   U96 : AOI22_X1 port map( A1 => c(14), A2 => n163, B1 => d(14), B2 => n160, 
                           ZN => n59);
   U97 : AOI22_X1 port map( A1 => c(15), A2 => n163, B1 => d(15), B2 => n160, 
                           ZN => n57);
   U98 : AOI22_X1 port map( A1 => c(16), A2 => n163, B1 => d(16), B2 => n160, 
                           ZN => n55);
   U99 : AOI22_X1 port map( A1 => c(17), A2 => n163, B1 => d(17), B2 => n160, 
                           ZN => n53);
   U100 : AOI22_X1 port map( A1 => c(18), A2 => n163, B1 => d(18), B2 => n160, 
                           ZN => n51);
   U101 : AOI22_X1 port map( A1 => c(19), A2 => n163, B1 => d(19), B2 => n160, 
                           ZN => n49);
   U102 : AOI22_X1 port map( A1 => c(20), A2 => n164, B1 => d(20), B2 => n161, 
                           ZN => n45);
   U103 : AOI22_X1 port map( A1 => c(21), A2 => n164, B1 => d(21), B2 => n161, 
                           ZN => n43);
   U104 : AOI22_X1 port map( A1 => c(22), A2 => n164, B1 => d(22), B2 => n161, 
                           ZN => n41);
   U105 : AOI22_X1 port map( A1 => c(23), A2 => n164, B1 => d(23), B2 => n161, 
                           ZN => n39);
   U106 : AOI22_X1 port map( A1 => c(24), A2 => n164, B1 => d(24), B2 => n161, 
                           ZN => n37);
   U107 : AOI22_X1 port map( A1 => c(25), A2 => n164, B1 => d(25), B2 => n161, 
                           ZN => n35);
   U108 : AOI22_X1 port map( A1 => c(26), A2 => n164, B1 => d(26), B2 => n161, 
                           ZN => n33);
   U109 : AOI22_X1 port map( A1 => c(27), A2 => n164, B1 => d(27), B2 => n161, 
                           ZN => n31);
   U110 : AOI22_X1 port map( A1 => c(28), A2 => n164, B1 => d(28), B2 => n161, 
                           ZN => n29);
   U111 : AOI22_X1 port map( A1 => c(29), A2 => n164, B1 => d(29), B2 => n161, 
                           ZN => n27);
   U112 : AOI22_X1 port map( A1 => c(30), A2 => n164, B1 => d(30), B2 => n161, 
                           ZN => n23);
   U113 : AOI22_X1 port map( A1 => c(31), A2 => n165, B1 => d(31), B2 => n162, 
                           ZN => n21);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_12 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_12;

architecture SYN_behavioral of reg_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n34, n35, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(0), QN => 
                           n36);
   U3 : BUF_X1 port map( A => n35, Z => n177);
   U4 : BUF_X1 port map( A => n35, Z => n176);
   U5 : BUF_X1 port map( A => n35, Z => n178);
   U6 : BUF_X1 port map( A => n34, Z => n179);
   U7 : BUF_X1 port map( A => n34, Z => n180);
   U8 : BUF_X1 port map( A => n34, Z => n181);
   U9 : NAND2_X1 port map( A1 => n182, A2 => n179, ZN => n35);
   U10 : OAI22_X1 port map( A1 => n181, A2 => n36, B1 => n178, B2 => n214, ZN 
                           => n99);
   U11 : INV_X1 port map( A => i(0), ZN => n214);
   U12 : OAI22_X1 port map( A1 => n181, A2 => n37, B1 => n178, B2 => n213, ZN 
                           => n98);
   U13 : INV_X1 port map( A => i(1), ZN => n213);
   U14 : OAI22_X1 port map( A1 => n181, A2 => n38, B1 => n178, B2 => n212, ZN 
                           => n97);
   U15 : INV_X1 port map( A => i(2), ZN => n212);
   U16 : OAI22_X1 port map( A1 => n181, A2 => n39, B1 => n178, B2 => n211, ZN 
                           => n96);
   U17 : INV_X1 port map( A => i(3), ZN => n211);
   U18 : OAI22_X1 port map( A1 => n181, A2 => n40, B1 => n178, B2 => n210, ZN 
                           => n95);
   U19 : INV_X1 port map( A => i(4), ZN => n210);
   U20 : OAI22_X1 port map( A1 => n181, A2 => n41, B1 => n178, B2 => n209, ZN 
                           => n94);
   U21 : INV_X1 port map( A => i(5), ZN => n209);
   U22 : OAI22_X1 port map( A1 => n181, A2 => n42, B1 => n178, B2 => n208, ZN 
                           => n93);
   U23 : INV_X1 port map( A => i(6), ZN => n208);
   U24 : OAI22_X1 port map( A1 => n180, A2 => n43, B1 => n178, B2 => n207, ZN 
                           => n92);
   U25 : INV_X1 port map( A => i(7), ZN => n207);
   U26 : OAI22_X1 port map( A1 => n180, A2 => n44, B1 => n177, B2 => n206, ZN 
                           => n91);
   U27 : INV_X1 port map( A => i(8), ZN => n206);
   U28 : OAI22_X1 port map( A1 => n180, A2 => n45, B1 => n177, B2 => n205, ZN 
                           => n90);
   U29 : INV_X1 port map( A => i(9), ZN => n205);
   U30 : OAI22_X1 port map( A1 => n180, A2 => n46, B1 => n177, B2 => n204, ZN 
                           => n89);
   U31 : INV_X1 port map( A => i(10), ZN => n204);
   U32 : OAI22_X1 port map( A1 => n180, A2 => n47, B1 => n177, B2 => n203, ZN 
                           => n88);
   U33 : INV_X1 port map( A => i(11), ZN => n203);
   U34 : OAI22_X1 port map( A1 => n180, A2 => n48, B1 => n177, B2 => n202, ZN 
                           => n87);
   U35 : INV_X1 port map( A => i(12), ZN => n202);
   U36 : OAI22_X1 port map( A1 => n180, A2 => n49, B1 => n177, B2 => n201, ZN 
                           => n86);
   U37 : INV_X1 port map( A => i(13), ZN => n201);
   U38 : OAI22_X1 port map( A1 => n180, A2 => n50, B1 => n177, B2 => n200, ZN 
                           => n85);
   U39 : INV_X1 port map( A => i(14), ZN => n200);
   U40 : OAI22_X1 port map( A1 => n180, A2 => n51, B1 => n177, B2 => n199, ZN 
                           => n84);
   U41 : INV_X1 port map( A => i(15), ZN => n199);
   U42 : OAI22_X1 port map( A1 => n180, A2 => n52, B1 => n177, B2 => n198, ZN 
                           => n83);
   U43 : INV_X1 port map( A => i(16), ZN => n198);
   U44 : OAI22_X1 port map( A1 => n180, A2 => n53, B1 => n177, B2 => n197, ZN 
                           => n82);
   U45 : INV_X1 port map( A => i(17), ZN => n197);
   U46 : OAI22_X1 port map( A1 => n180, A2 => n54, B1 => n177, B2 => n196, ZN 
                           => n81);
   U47 : INV_X1 port map( A => i(18), ZN => n196);
   U48 : OAI22_X1 port map( A1 => n180, A2 => n55, B1 => n177, B2 => n195, ZN 
                           => n80);
   U49 : INV_X1 port map( A => i(19), ZN => n195);
   U50 : OAI22_X1 port map( A1 => n179, A2 => n56, B1 => n176, B2 => n194, ZN 
                           => n79);
   U51 : INV_X1 port map( A => i(20), ZN => n194);
   U52 : OAI22_X1 port map( A1 => n179, A2 => n57, B1 => n176, B2 => n193, ZN 
                           => n78);
   U53 : INV_X1 port map( A => i(21), ZN => n193);
   U54 : OAI22_X1 port map( A1 => n179, A2 => n58, B1 => n176, B2 => n192, ZN 
                           => n77);
   U55 : INV_X1 port map( A => i(22), ZN => n192);
   U56 : OAI22_X1 port map( A1 => n179, A2 => n59, B1 => n176, B2 => n191, ZN 
                           => n76);
   U57 : INV_X1 port map( A => i(23), ZN => n191);
   U58 : OAI22_X1 port map( A1 => n179, A2 => n60, B1 => n176, B2 => n190, ZN 
                           => n75);
   U59 : INV_X1 port map( A => i(24), ZN => n190);
   U60 : OAI22_X1 port map( A1 => n179, A2 => n61, B1 => n176, B2 => n189, ZN 
                           => n74);
   U61 : INV_X1 port map( A => i(25), ZN => n189);
   U62 : OAI22_X1 port map( A1 => n179, A2 => n62, B1 => n176, B2 => n188, ZN 
                           => n73);
   U63 : INV_X1 port map( A => i(26), ZN => n188);
   U64 : OAI22_X1 port map( A1 => n179, A2 => n63, B1 => n176, B2 => n187, ZN 
                           => n72);
   U65 : INV_X1 port map( A => i(27), ZN => n187);
   U66 : OAI22_X1 port map( A1 => n179, A2 => n64, B1 => n176, B2 => n186, ZN 
                           => n71);
   U67 : INV_X1 port map( A => i(28), ZN => n186);
   U68 : OAI22_X1 port map( A1 => n179, A2 => n65, B1 => n176, B2 => n185, ZN 
                           => n70);
   U69 : INV_X1 port map( A => i(29), ZN => n185);
   U70 : OAI22_X1 port map( A1 => n179, A2 => n66, B1 => n176, B2 => n184, ZN 
                           => n69);
   U71 : INV_X1 port map( A => i(30), ZN => n184);
   U72 : OAI22_X1 port map( A1 => n179, A2 => n67, B1 => n176, B2 => n183, ZN 
                           => n68);
   U73 : INV_X1 port map( A => i(31), ZN => n183);
   U74 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n34);
   U75 : INV_X1 port map( A => reset, ZN => n182);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity reg_0 is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end reg_0;

architecture SYN_behavioral of reg_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n34, n35, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(31), QN =>
                           n67);
   temp_reg_30_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(30), QN =>
                           n66);
   temp_reg_29_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(29), QN =>
                           n65);
   temp_reg_28_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(28), QN =>
                           n64);
   temp_reg_27_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(27), QN =>
                           n63);
   temp_reg_26_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(26), QN =>
                           n62);
   temp_reg_25_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(25), QN =>
                           n61);
   temp_reg_24_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n97, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n98, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n99, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_3_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_1_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_8_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_9_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_0_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(0), QN => 
                           n36);
   temp_reg_5_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_6_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_7_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_4_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_2_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(2), QN => 
                           n38);
   U3 : BUF_X1 port map( A => n35, Z => n175);
   U4 : BUF_X1 port map( A => n35, Z => n174);
   U5 : BUF_X1 port map( A => n35, Z => n176);
   U6 : BUF_X1 port map( A => n34, Z => n178);
   U7 : BUF_X1 port map( A => n34, Z => n177);
   U8 : BUF_X1 port map( A => n34, Z => n179);
   U9 : NAND2_X1 port map( A1 => n180, A2 => n177, ZN => n35);
   U10 : INV_X1 port map( A => i(2), ZN => n190);
   U11 : OAI22_X1 port map( A1 => n179, A2 => n46, B1 => n176, B2 => n211, ZN 
                           => n99);
   U12 : INV_X1 port map( A => i(10), ZN => n211);
   U13 : OAI22_X1 port map( A1 => n179, A2 => n47, B1 => n176, B2 => n210, ZN 
                           => n98);
   U14 : INV_X1 port map( A => i(11), ZN => n210);
   U15 : OAI22_X1 port map( A1 => n179, A2 => n48, B1 => n176, B2 => n209, ZN 
                           => n97);
   U16 : INV_X1 port map( A => i(12), ZN => n209);
   U17 : OAI22_X1 port map( A1 => n179, A2 => n49, B1 => n176, B2 => n208, ZN 
                           => n96);
   U18 : INV_X1 port map( A => i(13), ZN => n208);
   U19 : OAI22_X1 port map( A1 => n179, A2 => n50, B1 => n176, B2 => n207, ZN 
                           => n95);
   U20 : INV_X1 port map( A => i(14), ZN => n207);
   U21 : OAI22_X1 port map( A1 => n179, A2 => n51, B1 => n176, B2 => n206, ZN 
                           => n94);
   U22 : INV_X1 port map( A => i(15), ZN => n206);
   U23 : OAI22_X1 port map( A1 => n179, A2 => n52, B1 => n176, B2 => n205, ZN 
                           => n93);
   U24 : INV_X1 port map( A => i(16), ZN => n205);
   U25 : OAI22_X1 port map( A1 => n178, A2 => n53, B1 => n176, B2 => n204, ZN 
                           => n92);
   U26 : INV_X1 port map( A => i(17), ZN => n204);
   U27 : OAI22_X1 port map( A1 => n177, A2 => n36, B1 => n174, B2 => n212, ZN 
                           => n77);
   U28 : INV_X1 port map( A => i(0), ZN => n212);
   U29 : OAI22_X1 port map( A1 => n177, A2 => n37, B1 => n174, B2 => n201, ZN 
                           => n76);
   U30 : INV_X1 port map( A => i(1), ZN => n201);
   U31 : OAI22_X1 port map( A1 => n177, A2 => n43, B1 => n174, B2 => n183, ZN 
                           => n70);
   U32 : INV_X1 port map( A => i(7), ZN => n183);
   U33 : OAI22_X1 port map( A1 => n177, A2 => n42, B1 => n174, B2 => n184, ZN 
                           => n71);
   U34 : INV_X1 port map( A => i(6), ZN => n184);
   U35 : OAI22_X1 port map( A1 => n177, A2 => n41, B1 => n174, B2 => n185, ZN 
                           => n72);
   U36 : INV_X1 port map( A => i(5), ZN => n185);
   U37 : OAI22_X1 port map( A1 => n177, A2 => n44, B1 => n174, B2 => n182, ZN 
                           => n69);
   U38 : INV_X1 port map( A => i(8), ZN => n182);
   U39 : OAI22_X1 port map( A1 => n177, A2 => n39, B1 => n174, B2 => n187, ZN 
                           => n74);
   U40 : INV_X1 port map( A => i(3), ZN => n187);
   U41 : OAI22_X1 port map( A1 => n177, A2 => n45, B1 => n174, B2 => n181, ZN 
                           => n68);
   U42 : INV_X1 port map( A => i(9), ZN => n181);
   U43 : OAI22_X1 port map( A1 => n177, A2 => n40, B1 => n174, B2 => n186, ZN 
                           => n73);
   U44 : INV_X1 port map( A => i(4), ZN => n186);
   U45 : OAI22_X1 port map( A1 => n178, A2 => n54, B1 => n175, B2 => n203, ZN 
                           => n91);
   U46 : INV_X1 port map( A => i(18), ZN => n203);
   U47 : OAI22_X1 port map( A1 => n178, A2 => n55, B1 => n175, B2 => n202, ZN 
                           => n90);
   U48 : INV_X1 port map( A => i(19), ZN => n202);
   U49 : OAI22_X1 port map( A1 => n178, A2 => n56, B1 => n175, B2 => n200, ZN 
                           => n89);
   U50 : INV_X1 port map( A => i(20), ZN => n200);
   U51 : OAI22_X1 port map( A1 => n178, A2 => n57, B1 => n175, B2 => n199, ZN 
                           => n88);
   U52 : INV_X1 port map( A => i(21), ZN => n199);
   U53 : OAI22_X1 port map( A1 => n178, A2 => n58, B1 => n175, B2 => n198, ZN 
                           => n87);
   U54 : INV_X1 port map( A => i(22), ZN => n198);
   U55 : OAI22_X1 port map( A1 => n178, A2 => n59, B1 => n175, B2 => n197, ZN 
                           => n86);
   U56 : INV_X1 port map( A => i(23), ZN => n197);
   U57 : OAI22_X1 port map( A1 => n178, A2 => n60, B1 => n175, B2 => n196, ZN 
                           => n85);
   U58 : INV_X1 port map( A => i(24), ZN => n196);
   U59 : OAI22_X1 port map( A1 => n178, A2 => n61, B1 => n175, B2 => n195, ZN 
                           => n84);
   U60 : INV_X1 port map( A => i(25), ZN => n195);
   U61 : OAI22_X1 port map( A1 => n178, A2 => n62, B1 => n175, B2 => n194, ZN 
                           => n83);
   U62 : INV_X1 port map( A => i(26), ZN => n194);
   U63 : OAI22_X1 port map( A1 => n178, A2 => n63, B1 => n175, B2 => n193, ZN 
                           => n82);
   U64 : INV_X1 port map( A => i(27), ZN => n193);
   U65 : OAI22_X1 port map( A1 => n178, A2 => n64, B1 => n175, B2 => n192, ZN 
                           => n81);
   U66 : INV_X1 port map( A => i(28), ZN => n192);
   U67 : OAI22_X1 port map( A1 => n178, A2 => n65, B1 => n175, B2 => n191, ZN 
                           => n80);
   U68 : INV_X1 port map( A => i(29), ZN => n191);
   U69 : OAI22_X1 port map( A1 => n177, A2 => n66, B1 => n174, B2 => n189, ZN 
                           => n79);
   U70 : INV_X1 port map( A => i(30), ZN => n189);
   U71 : OAI22_X1 port map( A1 => n177, A2 => n67, B1 => n174, B2 => n188, ZN 
                           => n78);
   U72 : INV_X1 port map( A => i(31), ZN => n188);
   U73 : OR2_X1 port map( A1 => load, A2 => reset, ZN => n34);
   U74 : OAI22_X1 port map( A1 => n177, A2 => n38, B1 => n174, B2 => n190, ZN 
                           => n75);
   U75 : INV_X1 port map( A => reset, ZN => n180);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity IR is

   port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 downto
         0);  o : out std_logic_vector (31 downto 0));

end IR;

architecture SYN_behavioral of IR is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n31, n32, n33, n34, n35, n97, n98, n99, n171, n172, n173
      , n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206 : std_logic;

begin
   
   temp_reg_31_inst : DFF_X1 port map( D => n68, CK => clock, Q => o(31), QN =>
                           n64);
   temp_reg_30_inst : DFF_X1 port map( D => n67, CK => clock, Q => o(30), QN =>
                           n97);
   temp_reg_29_inst : DFF_X1 port map( D => n69, CK => clock, Q => o(29), QN =>
                           n63);
   temp_reg_28_inst : DFF_X1 port map( D => n66, CK => clock, Q => o(28), QN =>
                           n98);
   temp_reg_27_inst : DFF_X1 port map( D => n70, CK => clock, Q => o(27), QN =>
                           n62);
   temp_reg_26_inst : DFF_X1 port map( D => n65, CK => clock, Q => o(26), QN =>
                           n99);
   temp_reg_24_inst : DFF_X1 port map( D => n72, CK => clock, Q => o(24), QN =>
                           n60);
   temp_reg_23_inst : DFF_X1 port map( D => n73, CK => clock, Q => o(23), QN =>
                           n59);
   temp_reg_22_inst : DFF_X1 port map( D => n74, CK => clock, Q => o(22), QN =>
                           n58);
   temp_reg_21_inst : DFF_X1 port map( D => n75, CK => clock, Q => o(21), QN =>
                           n57);
   temp_reg_20_inst : DFF_X1 port map( D => n76, CK => clock, Q => o(20), QN =>
                           n56);
   temp_reg_19_inst : DFF_X1 port map( D => n77, CK => clock, Q => o(19), QN =>
                           n55);
   temp_reg_18_inst : DFF_X1 port map( D => n78, CK => clock, Q => o(18), QN =>
                           n54);
   temp_reg_17_inst : DFF_X1 port map( D => n79, CK => clock, Q => o(17), QN =>
                           n53);
   temp_reg_16_inst : DFF_X1 port map( D => n80, CK => clock, Q => o(16), QN =>
                           n52);
   temp_reg_15_inst : DFF_X1 port map( D => n81, CK => clock, Q => o(15), QN =>
                           n51);
   temp_reg_14_inst : DFF_X1 port map( D => n82, CK => clock, Q => o(14), QN =>
                           n50);
   temp_reg_13_inst : DFF_X1 port map( D => n83, CK => clock, Q => o(13), QN =>
                           n49);
   temp_reg_12_inst : DFF_X1 port map( D => n84, CK => clock, Q => o(12), QN =>
                           n48);
   temp_reg_11_inst : DFF_X1 port map( D => n85, CK => clock, Q => o(11), QN =>
                           n47);
   temp_reg_10_inst : DFF_X1 port map( D => n86, CK => clock, Q => o(10), QN =>
                           n46);
   temp_reg_9_inst : DFF_X1 port map( D => n87, CK => clock, Q => o(9), QN => 
                           n45);
   temp_reg_8_inst : DFF_X1 port map( D => n88, CK => clock, Q => o(8), QN => 
                           n44);
   temp_reg_7_inst : DFF_X1 port map( D => n89, CK => clock, Q => o(7), QN => 
                           n43);
   temp_reg_6_inst : DFF_X1 port map( D => n90, CK => clock, Q => o(6), QN => 
                           n42);
   temp_reg_5_inst : DFF_X1 port map( D => n91, CK => clock, Q => o(5), QN => 
                           n41);
   temp_reg_4_inst : DFF_X1 port map( D => n92, CK => clock, Q => o(4), QN => 
                           n40);
   temp_reg_3_inst : DFF_X1 port map( D => n93, CK => clock, Q => o(3), QN => 
                           n39);
   temp_reg_2_inst : DFF_X1 port map( D => n94, CK => clock, Q => o(2), QN => 
                           n38);
   temp_reg_1_inst : DFF_X1 port map( D => n95, CK => clock, Q => o(1), QN => 
                           n37);
   temp_reg_0_inst : DFF_X1 port map( D => n96, CK => clock, Q => o(0), QN => 
                           n36);
   temp_reg_25_inst : DFF_X1 port map( D => n71, CK => clock, Q => o(25), QN =>
                           n61);
   U3 : BUF_X1 port map( A => n32, Z => n171);
   U4 : BUF_X1 port map( A => n32, Z => n172);
   U5 : BUF_X1 port map( A => n32, Z => n173);
   U6 : INV_X1 port map( A => reset, ZN => n177);
   U7 : NAND2_X1 port map( A1 => n177, A2 => n174, ZN => n32);
   U8 : BUF_X1 port map( A => n31, Z => n174);
   U9 : BUF_X1 port map( A => n31, Z => n175);
   U10 : BUF_X1 port map( A => n31, Z => n176);
   U11 : OAI22_X1 port map( A1 => n175, A2 => n36, B1 => n171, B2 => n206, ZN 
                           => n96);
   U12 : INV_X1 port map( A => i(0), ZN => n206);
   U13 : OAI22_X1 port map( A1 => n174, A2 => n37, B1 => n171, B2 => n205, ZN 
                           => n95);
   U14 : INV_X1 port map( A => i(1), ZN => n205);
   U15 : OAI22_X1 port map( A1 => n174, A2 => n38, B1 => n171, B2 => n204, ZN 
                           => n94);
   U16 : INV_X1 port map( A => i(2), ZN => n204);
   U17 : OAI22_X1 port map( A1 => n174, A2 => n39, B1 => n171, B2 => n203, ZN 
                           => n93);
   U18 : INV_X1 port map( A => i(3), ZN => n203);
   U19 : OAI22_X1 port map( A1 => n174, A2 => n40, B1 => n171, B2 => n202, ZN 
                           => n92);
   U20 : INV_X1 port map( A => i(4), ZN => n202);
   U21 : OAI22_X1 port map( A1 => n174, A2 => n41, B1 => n171, B2 => n201, ZN 
                           => n91);
   U22 : INV_X1 port map( A => i(5), ZN => n201);
   U23 : OAI22_X1 port map( A1 => n174, A2 => n42, B1 => n171, B2 => n200, ZN 
                           => n90);
   U24 : INV_X1 port map( A => i(6), ZN => n200);
   U25 : OAI22_X1 port map( A1 => n174, A2 => n43, B1 => n171, B2 => n199, ZN 
                           => n89);
   U26 : INV_X1 port map( A => i(7), ZN => n199);
   U27 : OAI22_X1 port map( A1 => n174, A2 => n44, B1 => n171, B2 => n198, ZN 
                           => n88);
   U28 : INV_X1 port map( A => i(8), ZN => n198);
   U29 : OAI22_X1 port map( A1 => n174, A2 => n45, B1 => n171, B2 => n197, ZN 
                           => n87);
   U30 : INV_X1 port map( A => i(9), ZN => n197);
   U31 : OAI22_X1 port map( A1 => n175, A2 => n46, B1 => n171, B2 => n196, ZN 
                           => n86);
   U32 : INV_X1 port map( A => i(10), ZN => n196);
   U33 : OAI22_X1 port map( A1 => n175, A2 => n47, B1 => n171, B2 => n195, ZN 
                           => n85);
   U34 : INV_X1 port map( A => i(11), ZN => n195);
   U35 : OAI22_X1 port map( A1 => n175, A2 => n48, B1 => n172, B2 => n194, ZN 
                           => n84);
   U36 : INV_X1 port map( A => i(12), ZN => n194);
   U37 : OAI22_X1 port map( A1 => n175, A2 => n49, B1 => n172, B2 => n193, ZN 
                           => n83);
   U38 : INV_X1 port map( A => i(13), ZN => n193);
   U39 : OAI22_X1 port map( A1 => n175, A2 => n50, B1 => n172, B2 => n192, ZN 
                           => n82);
   U40 : INV_X1 port map( A => i(14), ZN => n192);
   U41 : OAI22_X1 port map( A1 => n175, A2 => n51, B1 => n172, B2 => n191, ZN 
                           => n81);
   U42 : INV_X1 port map( A => i(15), ZN => n191);
   U43 : OAI22_X1 port map( A1 => n175, A2 => n52, B1 => n172, B2 => n190, ZN 
                           => n80);
   U44 : INV_X1 port map( A => i(16), ZN => n190);
   U45 : OAI22_X1 port map( A1 => n175, A2 => n53, B1 => n172, B2 => n189, ZN 
                           => n79);
   U46 : INV_X1 port map( A => i(17), ZN => n189);
   U47 : OAI22_X1 port map( A1 => n175, A2 => n54, B1 => n172, B2 => n188, ZN 
                           => n78);
   U48 : INV_X1 port map( A => i(18), ZN => n188);
   U49 : OAI22_X1 port map( A1 => n175, A2 => n55, B1 => n172, B2 => n187, ZN 
                           => n77);
   U50 : INV_X1 port map( A => i(19), ZN => n187);
   U51 : OAI22_X1 port map( A1 => n175, A2 => n56, B1 => n172, B2 => n186, ZN 
                           => n76);
   U52 : INV_X1 port map( A => i(20), ZN => n186);
   U53 : OAI22_X1 port map( A1 => n175, A2 => n57, B1 => n172, B2 => n185, ZN 
                           => n75);
   U54 : INV_X1 port map( A => i(21), ZN => n185);
   U55 : OAI22_X1 port map( A1 => n176, A2 => n58, B1 => n172, B2 => n184, ZN 
                           => n74);
   U56 : INV_X1 port map( A => i(22), ZN => n184);
   U57 : OAI22_X1 port map( A1 => n176, A2 => n59, B1 => n172, B2 => n183, ZN 
                           => n73);
   U58 : INV_X1 port map( A => i(23), ZN => n183);
   U59 : OAI22_X1 port map( A1 => n176, A2 => n61, B1 => n173, B2 => n181, ZN 
                           => n71);
   U60 : INV_X1 port map( A => i(25), ZN => n181);
   U61 : OAI22_X1 port map( A1 => n176, A2 => n60, B1 => n173, B2 => n182, ZN 
                           => n72);
   U62 : INV_X1 port map( A => i(24), ZN => n182);
   U63 : OAI22_X1 port map( A1 => n176, A2 => n62, B1 => n173, B2 => n180, ZN 
                           => n70);
   U64 : INV_X1 port map( A => i(27), ZN => n180);
   U65 : OAI22_X1 port map( A1 => n176, A2 => n63, B1 => n173, B2 => n179, ZN 
                           => n69);
   U66 : INV_X1 port map( A => i(29), ZN => n179);
   U67 : OAI22_X1 port map( A1 => n176, A2 => n64, B1 => n173, B2 => n178, ZN 
                           => n68);
   U68 : INV_X1 port map( A => i(31), ZN => n178);
   U69 : OAI211_X1 port map( C1 => n176, C2 => n99, A => n35, B => n177, ZN => 
                           n65);
   U70 : NAND2_X1 port map( A1 => i(26), A2 => n174, ZN => n35);
   U71 : OAI211_X1 port map( C1 => n176, C2 => n98, A => n34, B => n177, ZN => 
                           n66);
   U72 : NAND2_X1 port map( A1 => i(28), A2 => n174, ZN => n34);
   U73 : OAI211_X1 port map( C1 => n176, C2 => n97, A => n33, B => n177, ZN => 
                           n67);
   U74 : NAND2_X1 port map( A1 => i(30), A2 => n174, ZN => n33);
   U75 : OR2_X1 port map( A1 => reset, A2 => load, ZN => n31);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Mux21_0 is

   port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
         out std_logic_vector (31 downto 0));

end Mux21_0;

architecture SYN_Behavioral of Mux21_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n157, ZN => n145);
   U2 : CLKBUF_X1 port map( A => n158, Z => n156);
   U3 : CLKBUF_X1 port map( A => n158, Z => n155);
   U4 : INV_X1 port map( A => n157, ZN => n148);
   U5 : INV_X1 port map( A => n157, ZN => n147);
   U6 : BUF_X1 port map( A => n158, Z => n157);
   U7 : BUF_X1 port map( A => n158, Z => n154);
   U8 : BUF_X1 port map( A => n154, Z => n149);
   U9 : BUF_X1 port map( A => n158, Z => n153);
   U10 : BUF_X1 port map( A => n158, Z => n152);
   U11 : BUF_X1 port map( A => n153, Z => n151);
   U12 : BUF_X1 port map( A => n152, Z => n150);
   U13 : INV_X1 port map( A => n146, ZN => n158);
   U14 : BUF_X1 port map( A => sel, Z => n146);
   U15 : INV_X1 port map( A => n43, ZN => y(2));
   U16 : AOI22_X1 port map( A1 => a(2), A2 => n148, B1 => b(2), B2 => n151, ZN 
                           => n43);
   U17 : INV_X1 port map( A => n64, ZN => y(10));
   U18 : AOI22_X1 port map( A1 => a(10), A2 => n148, B1 => b(10), B2 => n156, 
                           ZN => n64);
   U19 : INV_X1 port map( A => n63, ZN => y(11));
   U20 : AOI22_X1 port map( A1 => a(11), A2 => n147, B1 => b(11), B2 => n156, 
                           ZN => n63);
   U21 : INV_X1 port map( A => n62, ZN => y(12));
   U22 : AOI22_X1 port map( A1 => a(12), A2 => n145, B1 => b(12), B2 => n156, 
                           ZN => n62);
   U23 : INV_X1 port map( A => n61, ZN => y(13));
   U24 : AOI22_X1 port map( A1 => a(13), A2 => n147, B1 => b(13), B2 => n155, 
                           ZN => n61);
   U25 : INV_X1 port map( A => n60, ZN => y(14));
   U26 : AOI22_X1 port map( A1 => a(14), A2 => n145, B1 => b(14), B2 => n155, 
                           ZN => n60);
   U27 : INV_X1 port map( A => n59, ZN => y(15));
   U28 : AOI22_X1 port map( A1 => a(15), A2 => n147, B1 => b(15), B2 => n155, 
                           ZN => n59);
   U29 : INV_X1 port map( A => n58, ZN => y(16));
   U30 : AOI22_X1 port map( A1 => a(16), A2 => n145, B1 => b(16), B2 => n155, 
                           ZN => n58);
   U31 : INV_X1 port map( A => n57, ZN => y(17));
   U32 : AOI22_X1 port map( A1 => a(17), A2 => n147, B1 => b(17), B2 => n154, 
                           ZN => n57);
   U33 : INV_X1 port map( A => n65, ZN => y(0));
   U34 : AOI22_X1 port map( A1 => a(0), A2 => n148, B1 => b(0), B2 => n156, ZN 
                           => n65);
   U35 : INV_X1 port map( A => n54, ZN => y(1));
   U36 : AOI22_X1 port map( A1 => a(1), A2 => n148, B1 => b(1), B2 => n154, ZN 
                           => n54);
   U37 : INV_X1 port map( A => n36, ZN => y(7));
   U38 : AOI22_X1 port map( A1 => a(7), A2 => n145, B1 => b(7), B2 => n149, ZN 
                           => n36);
   U39 : INV_X1 port map( A => n37, ZN => y(6));
   U40 : AOI22_X1 port map( A1 => a(6), A2 => n147, B1 => b(6), B2 => n149, ZN 
                           => n37);
   U41 : INV_X1 port map( A => n38, ZN => y(5));
   U42 : AOI22_X1 port map( A1 => a(5), A2 => n145, B1 => b(5), B2 => n150, ZN 
                           => n38);
   U43 : INV_X1 port map( A => n35, ZN => y(8));
   U44 : AOI22_X1 port map( A1 => a(8), A2 => n147, B1 => b(8), B2 => n149, ZN 
                           => n35);
   U45 : INV_X1 port map( A => n40, ZN => y(3));
   U46 : AOI22_X1 port map( A1 => a(3), A2 => n145, B1 => b(3), B2 => n150, ZN 
                           => n40);
   U47 : INV_X1 port map( A => n34, ZN => y(9));
   U48 : AOI22_X1 port map( A1 => n147, A2 => a(9), B1 => b(9), B2 => n149, ZN 
                           => n34);
   U49 : INV_X1 port map( A => n39, ZN => y(4));
   U50 : INV_X1 port map( A => n56, ZN => y(18));
   U51 : AOI22_X1 port map( A1 => a(18), A2 => n148, B1 => b(18), B2 => n154, 
                           ZN => n56);
   U52 : INV_X1 port map( A => n55, ZN => y(19));
   U53 : AOI22_X1 port map( A1 => a(19), A2 => n148, B1 => b(19), B2 => n154, 
                           ZN => n55);
   U54 : INV_X1 port map( A => n53, ZN => y(20));
   U55 : AOI22_X1 port map( A1 => a(20), A2 => n148, B1 => b(20), B2 => n153, 
                           ZN => n53);
   U56 : INV_X1 port map( A => n52, ZN => y(21));
   U57 : AOI22_X1 port map( A1 => a(21), A2 => n145, B1 => b(21), B2 => n153, 
                           ZN => n52);
   U58 : INV_X1 port map( A => n51, ZN => y(22));
   U59 : AOI22_X1 port map( A1 => a(22), A2 => n148, B1 => b(22), B2 => n153, 
                           ZN => n51);
   U60 : INV_X1 port map( A => n50, ZN => y(23));
   U61 : AOI22_X1 port map( A1 => a(23), A2 => n147, B1 => b(23), B2 => n153, 
                           ZN => n50);
   U62 : INV_X1 port map( A => n49, ZN => y(24));
   U63 : AOI22_X1 port map( A1 => a(24), A2 => n148, B1 => b(24), B2 => n152, 
                           ZN => n49);
   U64 : INV_X1 port map( A => n48, ZN => y(25));
   U65 : AOI22_X1 port map( A1 => a(25), A2 => n145, B1 => b(25), B2 => n152, 
                           ZN => n48);
   U66 : INV_X1 port map( A => n47, ZN => y(26));
   U67 : AOI22_X1 port map( A1 => a(26), A2 => n145, B1 => b(26), B2 => n152, 
                           ZN => n47);
   U68 : INV_X1 port map( A => n46, ZN => y(27));
   U69 : AOI22_X1 port map( A1 => a(27), A2 => n147, B1 => b(27), B2 => n152, 
                           ZN => n46);
   U70 : INV_X1 port map( A => n45, ZN => y(28));
   U71 : AOI22_X1 port map( A1 => a(28), A2 => n148, B1 => b(28), B2 => n151, 
                           ZN => n45);
   U72 : INV_X1 port map( A => n44, ZN => y(29));
   U73 : AOI22_X1 port map( A1 => a(29), A2 => n145, B1 => b(29), B2 => n151, 
                           ZN => n44);
   U74 : INV_X1 port map( A => n42, ZN => y(30));
   U75 : AOI22_X1 port map( A1 => a(30), A2 => n148, B1 => b(30), B2 => n151, 
                           ZN => n42);
   U76 : INV_X1 port map( A => n41, ZN => y(31));
   U77 : AOI22_X1 port map( A1 => a(31), A2 => n147, B1 => b(31), B2 => n150, 
                           ZN => n41);
   U78 : AOI22_X1 port map( A1 => a(4), A2 => n145, B1 => b(4), B2 => n150, ZN 
                           => n39);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Adder is

   port( A, B : in std_logic_vector (31 downto 0);  reset, Cin : in std_logic; 
         O : out std_logic_vector (31 downto 0);  Cout : out std_logic);

end Adder;

architecture SYN_Behavioral of Adder is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, O_0_port, N34
      , N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, 
      N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63
      , N64, N65, n7, n8, n9, n10, n_1351 : std_logic;

begin
   O <= ( O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, O_0_port );
   Cout <= O_31_port;
   
   add_1_root_add_26_2 : Adder_DW01_add_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), CI => Cin, SUM(31) => N65, 
                           SUM(30) => N64, SUM(29) => N63, SUM(28) => N62, 
                           SUM(27) => N61, SUM(26) => N60, SUM(25) => N59, 
                           SUM(24) => N58, SUM(23) => N57, SUM(22) => N56, 
                           SUM(21) => N55, SUM(20) => N54, SUM(19) => N53, 
                           SUM(18) => N52, SUM(17) => N51, SUM(16) => N50, 
                           SUM(15) => N49, SUM(14) => N48, SUM(13) => N47, 
                           SUM(12) => N46, SUM(11) => N45, SUM(10) => N44, 
                           SUM(9) => N43, SUM(8) => N42, SUM(7) => N41, SUM(6) 
                           => N40, SUM(5) => N39, SUM(4) => N38, SUM(3) => N37,
                           SUM(2) => N36, SUM(1) => N35, SUM(0) => N34, CO => 
                           n_1351);
   U2 : BUF_X1 port map( A => n10, Z => n7);
   U3 : BUF_X1 port map( A => n10, Z => n8);
   U4 : BUF_X1 port map( A => n10, Z => n9);
   U5 : AND2_X1 port map( A1 => N36, A2 => n8, ZN => O_2_port);
   U6 : AND2_X1 port map( A1 => N34, A2 => n7, ZN => O_0_port);
   U7 : AND2_X1 port map( A1 => N35, A2 => n7, ZN => O_1_port);
   U8 : AND2_X1 port map( A1 => N44, A2 => n7, ZN => O_10_port);
   U9 : AND2_X1 port map( A1 => N45, A2 => n7, ZN => O_11_port);
   U10 : AND2_X1 port map( A1 => N46, A2 => n7, ZN => O_12_port);
   U11 : AND2_X1 port map( A1 => N47, A2 => n7, ZN => O_13_port);
   U12 : AND2_X1 port map( A1 => N48, A2 => n7, ZN => O_14_port);
   U13 : AND2_X1 port map( A1 => N49, A2 => n7, ZN => O_15_port);
   U14 : AND2_X1 port map( A1 => N50, A2 => n7, ZN => O_16_port);
   U15 : AND2_X1 port map( A1 => N51, A2 => n7, ZN => O_17_port);
   U16 : AND2_X1 port map( A1 => N52, A2 => n7, ZN => O_18_port);
   U17 : AND2_X1 port map( A1 => N53, A2 => n7, ZN => O_19_port);
   U18 : AND2_X1 port map( A1 => N54, A2 => n8, ZN => O_20_port);
   U19 : AND2_X1 port map( A1 => N55, A2 => n8, ZN => O_21_port);
   U20 : AND2_X1 port map( A1 => N56, A2 => n8, ZN => O_22_port);
   U21 : AND2_X1 port map( A1 => N57, A2 => n8, ZN => O_23_port);
   U22 : AND2_X1 port map( A1 => N58, A2 => n8, ZN => O_24_port);
   U23 : AND2_X1 port map( A1 => N59, A2 => n8, ZN => O_25_port);
   U24 : AND2_X1 port map( A1 => N60, A2 => n8, ZN => O_26_port);
   U25 : AND2_X1 port map( A1 => N61, A2 => n8, ZN => O_27_port);
   U26 : AND2_X1 port map( A1 => N62, A2 => n8, ZN => O_28_port);
   U27 : AND2_X1 port map( A1 => N63, A2 => n8, ZN => O_29_port);
   U28 : AND2_X1 port map( A1 => N64, A2 => n8, ZN => O_30_port);
   U29 : AND2_X1 port map( A1 => N41, A2 => n9, ZN => O_7_port);
   U30 : AND2_X1 port map( A1 => N40, A2 => n9, ZN => O_6_port);
   U31 : AND2_X1 port map( A1 => N39, A2 => n9, ZN => O_5_port);
   U32 : AND2_X1 port map( A1 => N43, A2 => n9, ZN => O_9_port);
   U33 : AND2_X1 port map( A1 => N42, A2 => n9, ZN => O_8_port);
   U34 : AND2_X1 port map( A1 => N37, A2 => n9, ZN => O_3_port);
   U35 : AND2_X1 port map( A1 => N38, A2 => n9, ZN => O_4_port);
   U36 : INV_X1 port map( A => reset, ZN => n10);
   U37 : AND2_X1 port map( A1 => N65, A2 => n9, ZN => O_31_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity WBUnit is

   port( selwb : in std_logic;  ALUin, LOADDATA, AddressWfromMemory : in 
         std_logic_vector (31 downto 0);  MUXtoRF, AddressWtoDECODE : out 
         std_logic_vector (31 downto 0));

end WBUnit;

architecture SYN_structural of WBUnit is

   component Mux21_1
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;

begin
   AddressWtoDECODE <= ( AddressWfromMemory(31), AddressWfromMemory(30), 
      AddressWfromMemory(29), AddressWfromMemory(28), AddressWfromMemory(27), 
      AddressWfromMemory(26), AddressWfromMemory(25), AddressWfromMemory(24), 
      AddressWfromMemory(23), AddressWfromMemory(22), AddressWfromMemory(21), 
      AddressWfromMemory(20), AddressWfromMemory(19), AddressWfromMemory(18), 
      AddressWfromMemory(17), AddressWfromMemory(16), AddressWfromMemory(15), 
      AddressWfromMemory(14), AddressWfromMemory(13), AddressWfromMemory(12), 
      AddressWfromMemory(11), AddressWfromMemory(10), AddressWfromMemory(9), 
      AddressWfromMemory(8), AddressWfromMemory(7), AddressWfromMemory(6), 
      AddressWfromMemory(5), AddressWfromMemory(4), AddressWfromMemory(3), 
      AddressWfromMemory(2), AddressWfromMemory(1), AddressWfromMemory(0) );
   
   wbmux : Mux21_1 port map( a(31) => LOADDATA(31), a(30) => LOADDATA(30), 
                           a(29) => LOADDATA(29), a(28) => LOADDATA(28), a(27) 
                           => LOADDATA(27), a(26) => LOADDATA(26), a(25) => 
                           LOADDATA(25), a(24) => LOADDATA(24), a(23) => 
                           LOADDATA(23), a(22) => LOADDATA(22), a(21) => 
                           LOADDATA(21), a(20) => LOADDATA(20), a(19) => 
                           LOADDATA(19), a(18) => LOADDATA(18), a(17) => 
                           LOADDATA(17), a(16) => LOADDATA(16), a(15) => 
                           LOADDATA(15), a(14) => LOADDATA(14), a(13) => 
                           LOADDATA(13), a(12) => LOADDATA(12), a(11) => 
                           LOADDATA(11), a(10) => LOADDATA(10), a(9) => 
                           LOADDATA(9), a(8) => LOADDATA(8), a(7) => 
                           LOADDATA(7), a(6) => LOADDATA(6), a(5) => 
                           LOADDATA(5), a(4) => LOADDATA(4), a(3) => 
                           LOADDATA(3), a(2) => LOADDATA(2), a(1) => 
                           LOADDATA(1), a(0) => LOADDATA(0), b(31) => ALUin(31)
                           , b(30) => ALUin(30), b(29) => ALUin(29), b(28) => 
                           ALUin(28), b(27) => ALUin(27), b(26) => ALUin(26), 
                           b(25) => ALUin(25), b(24) => ALUin(24), b(23) => 
                           ALUin(23), b(22) => ALUin(22), b(21) => ALUin(21), 
                           b(20) => ALUin(20), b(19) => ALUin(19), b(18) => 
                           ALUin(18), b(17) => ALUin(17), b(16) => ALUin(16), 
                           b(15) => ALUin(15), b(14) => ALUin(14), b(13) => 
                           ALUin(13), b(12) => ALUin(12), b(11) => ALUin(11), 
                           b(10) => ALUin(10), b(9) => ALUin(9), b(8) => 
                           ALUin(8), b(7) => ALUin(7), b(6) => ALUin(6), b(5) 
                           => ALUin(5), b(4) => ALUin(4), b(3) => ALUin(3), 
                           b(2) => ALUin(2), b(1) => ALUin(1), b(0) => ALUin(0)
                           , sel => selwb, y(31) => MUXtoRF(31), y(30) => 
                           MUXtoRF(30), y(29) => MUXtoRF(29), y(28) => 
                           MUXtoRF(28), y(27) => MUXtoRF(27), y(26) => 
                           MUXtoRF(26), y(25) => MUXtoRF(25), y(24) => 
                           MUXtoRF(24), y(23) => MUXtoRF(23), y(22) => 
                           MUXtoRF(22), y(21) => MUXtoRF(21), y(20) => 
                           MUXtoRF(20), y(19) => MUXtoRF(19), y(18) => 
                           MUXtoRF(18), y(17) => MUXtoRF(17), y(16) => 
                           MUXtoRF(16), y(15) => MUXtoRF(15), y(14) => 
                           MUXtoRF(14), y(13) => MUXtoRF(13), y(12) => 
                           MUXtoRF(12), y(11) => MUXtoRF(11), y(10) => 
                           MUXtoRF(10), y(9) => MUXtoRF(9), y(8) => MUXtoRF(8),
                           y(7) => MUXtoRF(7), y(6) => MUXtoRF(6), y(5) => 
                           MUXtoRF(5), y(4) => MUXtoRF(4), y(3) => MUXtoRF(3), 
                           y(2) => MUXtoRF(2), y(1) => MUXtoRF(1), y(0) => 
                           MUXtoRF(0));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity memoryUnit is

   port( clock, reset, en4 : in std_logic;  ALUout, DRAMout, 
         AddressWfromEXECUTE : in std_logic_vector (31 downto 0);  LOADDATA, 
         ALUtoWBMUX, AddressWtoWB : out std_logic_vector (31 downto 0));

end memoryUnit;

architecture SYN_structural of memoryUnit is

   component reg_1
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_2
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_3
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;

begin
   
   LMD_REG : reg_3 port map( clock => clock, reset => reset, load => en4, i(31)
                           => DRAMout(31), i(30) => DRAMout(30), i(29) => 
                           DRAMout(29), i(28) => DRAMout(28), i(27) => 
                           DRAMout(27), i(26) => DRAMout(26), i(25) => 
                           DRAMout(25), i(24) => DRAMout(24), i(23) => 
                           DRAMout(23), i(22) => DRAMout(22), i(21) => 
                           DRAMout(21), i(20) => DRAMout(20), i(19) => 
                           DRAMout(19), i(18) => DRAMout(18), i(17) => 
                           DRAMout(17), i(16) => DRAMout(16), i(15) => 
                           DRAMout(15), i(14) => DRAMout(14), i(13) => 
                           DRAMout(13), i(12) => DRAMout(12), i(11) => 
                           DRAMout(11), i(10) => DRAMout(10), i(9) => 
                           DRAMout(9), i(8) => DRAMout(8), i(7) => DRAMout(7), 
                           i(6) => DRAMout(6), i(5) => DRAMout(5), i(4) => 
                           DRAMout(4), i(3) => DRAMout(3), i(2) => DRAMout(2), 
                           i(1) => DRAMout(1), i(0) => DRAMout(0), o(31) => 
                           LOADDATA(31), o(30) => LOADDATA(30), o(29) => 
                           LOADDATA(29), o(28) => LOADDATA(28), o(27) => 
                           LOADDATA(27), o(26) => LOADDATA(26), o(25) => 
                           LOADDATA(25), o(24) => LOADDATA(24), o(23) => 
                           LOADDATA(23), o(22) => LOADDATA(22), o(21) => 
                           LOADDATA(21), o(20) => LOADDATA(20), o(19) => 
                           LOADDATA(19), o(18) => LOADDATA(18), o(17) => 
                           LOADDATA(17), o(16) => LOADDATA(16), o(15) => 
                           LOADDATA(15), o(14) => LOADDATA(14), o(13) => 
                           LOADDATA(13), o(12) => LOADDATA(12), o(11) => 
                           LOADDATA(11), o(10) => LOADDATA(10), o(9) => 
                           LOADDATA(9), o(8) => LOADDATA(8), o(7) => 
                           LOADDATA(7), o(6) => LOADDATA(6), o(5) => 
                           LOADDATA(5), o(4) => LOADDATA(4), o(3) => 
                           LOADDATA(3), o(2) => LOADDATA(2), o(1) => 
                           LOADDATA(1), o(0) => LOADDATA(0));
   ALUout_REG : reg_2 port map( clock => clock, reset => reset, load => en4, 
                           i(31) => ALUout(31), i(30) => ALUout(30), i(29) => 
                           ALUout(29), i(28) => ALUout(28), i(27) => ALUout(27)
                           , i(26) => ALUout(26), i(25) => ALUout(25), i(24) =>
                           ALUout(24), i(23) => ALUout(23), i(22) => ALUout(22)
                           , i(21) => ALUout(21), i(20) => ALUout(20), i(19) =>
                           ALUout(19), i(18) => ALUout(18), i(17) => ALUout(17)
                           , i(16) => ALUout(16), i(15) => ALUout(15), i(14) =>
                           ALUout(14), i(13) => ALUout(13), i(12) => ALUout(12)
                           , i(11) => ALUout(11), i(10) => ALUout(10), i(9) => 
                           ALUout(9), i(8) => ALUout(8), i(7) => ALUout(7), 
                           i(6) => ALUout(6), i(5) => ALUout(5), i(4) => 
                           ALUout(4), i(3) => ALUout(3), i(2) => ALUout(2), 
                           i(1) => ALUout(1), i(0) => ALUout(0), o(31) => 
                           ALUtoWBMUX(31), o(30) => ALUtoWBMUX(30), o(29) => 
                           ALUtoWBMUX(29), o(28) => ALUtoWBMUX(28), o(27) => 
                           ALUtoWBMUX(27), o(26) => ALUtoWBMUX(26), o(25) => 
                           ALUtoWBMUX(25), o(24) => ALUtoWBMUX(24), o(23) => 
                           ALUtoWBMUX(23), o(22) => ALUtoWBMUX(22), o(21) => 
                           ALUtoWBMUX(21), o(20) => ALUtoWBMUX(20), o(19) => 
                           ALUtoWBMUX(19), o(18) => ALUtoWBMUX(18), o(17) => 
                           ALUtoWBMUX(17), o(16) => ALUtoWBMUX(16), o(15) => 
                           ALUtoWBMUX(15), o(14) => ALUtoWBMUX(14), o(13) => 
                           ALUtoWBMUX(13), o(12) => ALUtoWBMUX(12), o(11) => 
                           ALUtoWBMUX(11), o(10) => ALUtoWBMUX(10), o(9) => 
                           ALUtoWBMUX(9), o(8) => ALUtoWBMUX(8), o(7) => 
                           ALUtoWBMUX(7), o(6) => ALUtoWBMUX(6), o(5) => 
                           ALUtoWBMUX(5), o(4) => ALUtoWBMUX(4), o(3) => 
                           ALUtoWBMUX(3), o(2) => ALUtoWBMUX(2), o(1) => 
                           ALUtoWBMUX(1), o(0) => ALUtoWBMUX(0));
   AddressW_REG : reg_1 port map( clock => clock, reset => reset, load => en4, 
                           i(31) => AddressWfromEXECUTE(31), i(30) => 
                           AddressWfromEXECUTE(30), i(29) => 
                           AddressWfromEXECUTE(29), i(28) => 
                           AddressWfromEXECUTE(28), i(27) => 
                           AddressWfromEXECUTE(27), i(26) => 
                           AddressWfromEXECUTE(26), i(25) => 
                           AddressWfromEXECUTE(25), i(24) => 
                           AddressWfromEXECUTE(24), i(23) => 
                           AddressWfromEXECUTE(23), i(22) => 
                           AddressWfromEXECUTE(22), i(21) => 
                           AddressWfromEXECUTE(21), i(20) => 
                           AddressWfromEXECUTE(20), i(19) => 
                           AddressWfromEXECUTE(19), i(18) => 
                           AddressWfromEXECUTE(18), i(17) => 
                           AddressWfromEXECUTE(17), i(16) => 
                           AddressWfromEXECUTE(16), i(15) => 
                           AddressWfromEXECUTE(15), i(14) => 
                           AddressWfromEXECUTE(14), i(13) => 
                           AddressWfromEXECUTE(13), i(12) => 
                           AddressWfromEXECUTE(12), i(11) => 
                           AddressWfromEXECUTE(11), i(10) => 
                           AddressWfromEXECUTE(10), i(9) => 
                           AddressWfromEXECUTE(9), i(8) => 
                           AddressWfromEXECUTE(8), i(7) => 
                           AddressWfromEXECUTE(7), i(6) => 
                           AddressWfromEXECUTE(6), i(5) => 
                           AddressWfromEXECUTE(5), i(4) => 
                           AddressWfromEXECUTE(4), i(3) => 
                           AddressWfromEXECUTE(3), i(2) => 
                           AddressWfromEXECUTE(2), i(1) => 
                           AddressWfromEXECUTE(1), i(0) => 
                           AddressWfromEXECUTE(0), o(31) => AddressWtoWB(31), 
                           o(30) => AddressWtoWB(30), o(29) => AddressWtoWB(29)
                           , o(28) => AddressWtoWB(28), o(27) => 
                           AddressWtoWB(27), o(26) => AddressWtoWB(26), o(25) 
                           => AddressWtoWB(25), o(24) => AddressWtoWB(24), 
                           o(23) => AddressWtoWB(23), o(22) => AddressWtoWB(22)
                           , o(21) => AddressWtoWB(21), o(20) => 
                           AddressWtoWB(20), o(19) => AddressWtoWB(19), o(18) 
                           => AddressWtoWB(18), o(17) => AddressWtoWB(17), 
                           o(16) => AddressWtoWB(16), o(15) => AddressWtoWB(15)
                           , o(14) => AddressWtoWB(14), o(13) => 
                           AddressWtoWB(13), o(12) => AddressWtoWB(12), o(11) 
                           => AddressWtoWB(11), o(10) => AddressWtoWB(10), o(9)
                           => AddressWtoWB(9), o(8) => AddressWtoWB(8), o(7) =>
                           AddressWtoWB(7), o(6) => AddressWtoWB(6), o(5) => 
                           AddressWtoWB(5), o(4) => AddressWtoWB(4), o(3) => 
                           AddressWtoWB(3), o(2) => AddressWtoWB(2), o(1) => 
                           AddressWtoWB(1), o(0) => AddressWtoWB(0));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity executeUnit_M32_C4 is

   port( clock, reset, en3, Mux1Sel, Mux2Sel : in std_logic;  ALUCODE : in 
         std_logic_vector (3 downto 0);  OUT1RF, OUT2RF, IMMEDIATE, 
         NPCFromDecode, AddressWfromDecode : in std_logic_vector (31 downto 0);
         ALUtoMEMORY, OUT2RFtoMEMORY, AddressWtoMEMORY : out std_logic_vector 
         (31 downto 0));

end executeUnit_M32_C4;

architecture SYN_structural of executeUnit_M32_C4 is

   component reg_4
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_5
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_6
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component ALU_M32_C4
      port( CODE : in std_logic_vector (3 downto 0);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Mux21_2
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component Mux21_3
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component Mux21_4
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal X_Logic0_port, MUX2out_31_port, MUX2out_30_port, MUX2out_29_port, 
      MUX2out_28_port, MUX2out_27_port, MUX2out_26_port, MUX2out_25_port, 
      MUX2out_24_port, MUX2out_23_port, MUX2out_22_port, MUX2out_21_port, 
      MUX2out_20_port, MUX2out_19_port, MUX2out_18_port, MUX2out_17_port, 
      MUX2out_16_port, MUX2out_15_port, MUX2out_14_port, MUX2out_13_port, 
      MUX2out_12_port, MUX2out_11_port, MUX2out_10_port, MUX2out_9_port, 
      MUX2out_8_port, MUX2out_7_port, MUX2out_6_port, MUX2out_5_port, 
      MUX2out_4_port, MUX2out_3_port, MUX2out_2_port, MUX2out_1_port, 
      MUX2out_0_port, MUXNPCout_31_port, MUXNPCout_30_port, MUXNPCout_29_port, 
      MUXNPCout_28_port, MUXNPCout_27_port, MUXNPCout_26_port, 
      MUXNPCout_25_port, MUXNPCout_24_port, MUXNPCout_23_port, 
      MUXNPCout_22_port, MUXNPCout_21_port, MUXNPCout_20_port, 
      MUXNPCout_19_port, MUXNPCout_18_port, MUXNPCout_17_port, 
      MUXNPCout_16_port, MUXNPCout_15_port, MUXNPCout_14_port, 
      MUXNPCout_13_port, MUXNPCout_12_port, MUXNPCout_11_port, 
      MUXNPCout_10_port, MUXNPCout_9_port, MUXNPCout_8_port, MUXNPCout_7_port, 
      MUXNPCout_6_port, MUXNPCout_5_port, MUXNPCout_4_port, MUXNPCout_3_port, 
      MUXNPCout_2_port, MUXNPCout_1_port, MUXNPCout_0_port, MUXWITH4out_31_port
      , MUXWITH4out_30_port, MUXWITH4out_29_port, MUXWITH4out_28_port, 
      MUXWITH4out_27_port, MUXWITH4out_26_port, MUXWITH4out_25_port, 
      MUXWITH4out_24_port, MUXWITH4out_23_port, MUXWITH4out_22_port, 
      MUXWITH4out_21_port, MUXWITH4out_20_port, MUXWITH4out_19_port, 
      MUXWITH4out_18_port, MUXWITH4out_17_port, MUXWITH4out_16_port, 
      MUXWITH4out_15_port, MUXWITH4out_14_port, MUXWITH4out_13_port, 
      MUXWITH4out_12_port, MUXWITH4out_11_port, MUXWITH4out_10_port, 
      MUXWITH4out_9_port, MUXWITH4out_8_port, MUXWITH4out_7_port, 
      MUXWITH4out_6_port, MUXWITH4out_5_port, MUXWITH4out_4_port, 
      MUXWITH4out_3_port, MUXWITH4out_2_port, MUXWITH4out_1_port, 
      MUXWITH4out_0_port, ALUout_31_port, ALUout_30_port, ALUout_29_port, 
      ALUout_28_port, ALUout_27_port, ALUout_26_port, ALUout_25_port, 
      ALUout_24_port, ALUout_23_port, ALUout_22_port, ALUout_21_port, 
      ALUout_20_port, ALUout_19_port, ALUout_18_port, ALUout_17_port, 
      ALUout_16_port, ALUout_15_port, ALUout_14_port, ALUout_13_port, 
      ALUout_12_port, ALUout_11_port, ALUout_10_port, ALUout_9_port, 
      ALUout_8_port, ALUout_7_port, ALUout_6_port, ALUout_5_port, ALUout_4_port
      , ALUout_3_port, ALUout_2_port, ALUout_1_port, ALUout_0_port : std_logic;

begin
   
   X_Logic0_port <= '0';
   MUX : Mux21_4 port map( a(31) => OUT2RF(31), a(30) => OUT2RF(30), a(29) => 
                           OUT2RF(29), a(28) => OUT2RF(28), a(27) => OUT2RF(27)
                           , a(26) => OUT2RF(26), a(25) => OUT2RF(25), a(24) =>
                           OUT2RF(24), a(23) => OUT2RF(23), a(22) => OUT2RF(22)
                           , a(21) => OUT2RF(21), a(20) => OUT2RF(20), a(19) =>
                           OUT2RF(19), a(18) => OUT2RF(18), a(17) => OUT2RF(17)
                           , a(16) => OUT2RF(16), a(15) => OUT2RF(15), a(14) =>
                           OUT2RF(14), a(13) => OUT2RF(13), a(12) => OUT2RF(12)
                           , a(11) => OUT2RF(11), a(10) => OUT2RF(10), a(9) => 
                           OUT2RF(9), a(8) => OUT2RF(8), a(7) => OUT2RF(7), 
                           a(6) => OUT2RF(6), a(5) => OUT2RF(5), a(4) => 
                           OUT2RF(4), a(3) => OUT2RF(3), a(2) => OUT2RF(2), 
                           a(1) => OUT2RF(1), a(0) => OUT2RF(0), b(31) => 
                           IMMEDIATE(31), b(30) => IMMEDIATE(30), b(29) => 
                           IMMEDIATE(29), b(28) => IMMEDIATE(28), b(27) => 
                           IMMEDIATE(27), b(26) => IMMEDIATE(26), b(25) => 
                           IMMEDIATE(25), b(24) => IMMEDIATE(24), b(23) => 
                           IMMEDIATE(23), b(22) => IMMEDIATE(22), b(21) => 
                           IMMEDIATE(21), b(20) => IMMEDIATE(20), b(19) => 
                           IMMEDIATE(19), b(18) => IMMEDIATE(18), b(17) => 
                           IMMEDIATE(17), b(16) => IMMEDIATE(16), b(15) => 
                           IMMEDIATE(15), b(14) => IMMEDIATE(14), b(13) => 
                           IMMEDIATE(13), b(12) => IMMEDIATE(12), b(11) => 
                           IMMEDIATE(11), b(10) => IMMEDIATE(10), b(9) => 
                           IMMEDIATE(9), b(8) => IMMEDIATE(8), b(7) => 
                           IMMEDIATE(7), b(6) => IMMEDIATE(6), b(5) => 
                           IMMEDIATE(5), b(4) => IMMEDIATE(4), b(3) => 
                           IMMEDIATE(3), b(2) => IMMEDIATE(2), b(1) => 
                           IMMEDIATE(1), b(0) => IMMEDIATE(0), sel => Mux2Sel, 
                           y(31) => MUX2out_31_port, y(30) => MUX2out_30_port, 
                           y(29) => MUX2out_29_port, y(28) => MUX2out_28_port, 
                           y(27) => MUX2out_27_port, y(26) => MUX2out_26_port, 
                           y(25) => MUX2out_25_port, y(24) => MUX2out_24_port, 
                           y(23) => MUX2out_23_port, y(22) => MUX2out_22_port, 
                           y(21) => MUX2out_21_port, y(20) => MUX2out_20_port, 
                           y(19) => MUX2out_19_port, y(18) => MUX2out_18_port, 
                           y(17) => MUX2out_17_port, y(16) => MUX2out_16_port, 
                           y(15) => MUX2out_15_port, y(14) => MUX2out_14_port, 
                           y(13) => MUX2out_13_port, y(12) => MUX2out_12_port, 
                           y(11) => MUX2out_11_port, y(10) => MUX2out_10_port, 
                           y(9) => MUX2out_9_port, y(8) => MUX2out_8_port, y(7)
                           => MUX2out_7_port, y(6) => MUX2out_6_port, y(5) => 
                           MUX2out_5_port, y(4) => MUX2out_4_port, y(3) => 
                           MUX2out_3_port, y(2) => MUX2out_2_port, y(1) => 
                           MUX2out_1_port, y(0) => MUX2out_0_port);
   MUXNPC : Mux21_3 port map( a(31) => NPCFromDecode(31), a(30) => 
                           NPCFromDecode(30), a(29) => NPCFromDecode(29), a(28)
                           => NPCFromDecode(28), a(27) => NPCFromDecode(27), 
                           a(26) => NPCFromDecode(26), a(25) => 
                           NPCFromDecode(25), a(24) => NPCFromDecode(24), a(23)
                           => NPCFromDecode(23), a(22) => NPCFromDecode(22), 
                           a(21) => NPCFromDecode(21), a(20) => 
                           NPCFromDecode(20), a(19) => NPCFromDecode(19), a(18)
                           => NPCFromDecode(18), a(17) => NPCFromDecode(17), 
                           a(16) => NPCFromDecode(16), a(15) => 
                           NPCFromDecode(15), a(14) => NPCFromDecode(14), a(13)
                           => NPCFromDecode(13), a(12) => NPCFromDecode(12), 
                           a(11) => NPCFromDecode(11), a(10) => 
                           NPCFromDecode(10), a(9) => NPCFromDecode(9), a(8) =>
                           NPCFromDecode(8), a(7) => NPCFromDecode(7), a(6) => 
                           NPCFromDecode(6), a(5) => NPCFromDecode(5), a(4) => 
                           NPCFromDecode(4), a(3) => NPCFromDecode(3), a(2) => 
                           NPCFromDecode(2), a(1) => NPCFromDecode(1), a(0) => 
                           NPCFromDecode(0), b(31) => OUT1RF(31), b(30) => 
                           OUT1RF(30), b(29) => OUT1RF(29), b(28) => OUT1RF(28)
                           , b(27) => OUT1RF(27), b(26) => OUT1RF(26), b(25) =>
                           OUT1RF(25), b(24) => OUT1RF(24), b(23) => OUT1RF(23)
                           , b(22) => OUT1RF(22), b(21) => OUT1RF(21), b(20) =>
                           OUT1RF(20), b(19) => OUT1RF(19), b(18) => OUT1RF(18)
                           , b(17) => OUT1RF(17), b(16) => OUT1RF(16), b(15) =>
                           OUT1RF(15), b(14) => OUT1RF(14), b(13) => OUT1RF(13)
                           , b(12) => OUT1RF(12), b(11) => OUT1RF(11), b(10) =>
                           OUT1RF(10), b(9) => OUT1RF(9), b(8) => OUT1RF(8), 
                           b(7) => OUT1RF(7), b(6) => OUT1RF(6), b(5) => 
                           OUT1RF(5), b(4) => OUT1RF(4), b(3) => OUT1RF(3), 
                           b(2) => OUT1RF(2), b(1) => OUT1RF(1), b(0) => 
                           OUT1RF(0), sel => Mux1Sel, y(31) => 
                           MUXNPCout_31_port, y(30) => MUXNPCout_30_port, y(29)
                           => MUXNPCout_29_port, y(28) => MUXNPCout_28_port, 
                           y(27) => MUXNPCout_27_port, y(26) => 
                           MUXNPCout_26_port, y(25) => MUXNPCout_25_port, y(24)
                           => MUXNPCout_24_port, y(23) => MUXNPCout_23_port, 
                           y(22) => MUXNPCout_22_port, y(21) => 
                           MUXNPCout_21_port, y(20) => MUXNPCout_20_port, y(19)
                           => MUXNPCout_19_port, y(18) => MUXNPCout_18_port, 
                           y(17) => MUXNPCout_17_port, y(16) => 
                           MUXNPCout_16_port, y(15) => MUXNPCout_15_port, y(14)
                           => MUXNPCout_14_port, y(13) => MUXNPCout_13_port, 
                           y(12) => MUXNPCout_12_port, y(11) => 
                           MUXNPCout_11_port, y(10) => MUXNPCout_10_port, y(9) 
                           => MUXNPCout_9_port, y(8) => MUXNPCout_8_port, y(7) 
                           => MUXNPCout_7_port, y(6) => MUXNPCout_6_port, y(5) 
                           => MUXNPCout_5_port, y(4) => MUXNPCout_4_port, y(3) 
                           => MUXNPCout_3_port, y(2) => MUXNPCout_2_port, y(1) 
                           => MUXNPCout_1_port, y(0) => MUXNPCout_0_port);
   MUXWITH4 : Mux21_2 port map( a(31) => X_Logic0_port, a(30) => X_Logic0_port,
                           a(29) => X_Logic0_port, a(28) => X_Logic0_port, 
                           a(27) => X_Logic0_port, a(26) => X_Logic0_port, 
                           a(25) => X_Logic0_port, a(24) => X_Logic0_port, 
                           a(23) => X_Logic0_port, a(22) => X_Logic0_port, 
                           a(21) => X_Logic0_port, a(20) => X_Logic0_port, 
                           a(19) => X_Logic0_port, a(18) => X_Logic0_port, 
                           a(17) => X_Logic0_port, a(16) => X_Logic0_port, 
                           a(15) => X_Logic0_port, a(14) => X_Logic0_port, 
                           a(13) => X_Logic0_port, a(12) => X_Logic0_port, 
                           a(11) => X_Logic0_port, a(10) => X_Logic0_port, a(9)
                           => X_Logic0_port, a(8) => X_Logic0_port, a(7) => 
                           X_Logic0_port, a(6) => X_Logic0_port, a(5) => 
                           X_Logic0_port, a(4) => X_Logic0_port, a(3) => 
                           X_Logic0_port, a(2) => X_Logic0_port, a(1) => 
                           X_Logic0_port, a(0) => X_Logic0_port, b(31) => 
                           MUX2out_31_port, b(30) => MUX2out_30_port, b(29) => 
                           MUX2out_29_port, b(28) => MUX2out_28_port, b(27) => 
                           MUX2out_27_port, b(26) => MUX2out_26_port, b(25) => 
                           MUX2out_25_port, b(24) => MUX2out_24_port, b(23) => 
                           MUX2out_23_port, b(22) => MUX2out_22_port, b(21) => 
                           MUX2out_21_port, b(20) => MUX2out_20_port, b(19) => 
                           MUX2out_19_port, b(18) => MUX2out_18_port, b(17) => 
                           MUX2out_17_port, b(16) => MUX2out_16_port, b(15) => 
                           MUX2out_15_port, b(14) => MUX2out_14_port, b(13) => 
                           MUX2out_13_port, b(12) => MUX2out_12_port, b(11) => 
                           MUX2out_11_port, b(10) => MUX2out_10_port, b(9) => 
                           MUX2out_9_port, b(8) => MUX2out_8_port, b(7) => 
                           MUX2out_7_port, b(6) => MUX2out_6_port, b(5) => 
                           MUX2out_5_port, b(4) => MUX2out_4_port, b(3) => 
                           MUX2out_3_port, b(2) => MUX2out_2_port, b(1) => 
                           MUX2out_1_port, b(0) => MUX2out_0_port, sel => 
                           Mux1Sel, y(31) => MUXWITH4out_31_port, y(30) => 
                           MUXWITH4out_30_port, y(29) => MUXWITH4out_29_port, 
                           y(28) => MUXWITH4out_28_port, y(27) => 
                           MUXWITH4out_27_port, y(26) => MUXWITH4out_26_port, 
                           y(25) => MUXWITH4out_25_port, y(24) => 
                           MUXWITH4out_24_port, y(23) => MUXWITH4out_23_port, 
                           y(22) => MUXWITH4out_22_port, y(21) => 
                           MUXWITH4out_21_port, y(20) => MUXWITH4out_20_port, 
                           y(19) => MUXWITH4out_19_port, y(18) => 
                           MUXWITH4out_18_port, y(17) => MUXWITH4out_17_port, 
                           y(16) => MUXWITH4out_16_port, y(15) => 
                           MUXWITH4out_15_port, y(14) => MUXWITH4out_14_port, 
                           y(13) => MUXWITH4out_13_port, y(12) => 
                           MUXWITH4out_12_port, y(11) => MUXWITH4out_11_port, 
                           y(10) => MUXWITH4out_10_port, y(9) => 
                           MUXWITH4out_9_port, y(8) => MUXWITH4out_8_port, y(7)
                           => MUXWITH4out_7_port, y(6) => MUXWITH4out_6_port, 
                           y(5) => MUXWITH4out_5_port, y(4) => 
                           MUXWITH4out_4_port, y(3) => MUXWITH4out_3_port, y(2)
                           => MUXWITH4out_2_port, y(1) => MUXWITH4out_1_port, 
                           y(0) => MUXWITH4out_0_port);
   ALUset : ALU_M32_C4 port map( CODE(3) => ALUCODE(3), CODE(2) => ALUCODE(2), 
                           CODE(1) => ALUCODE(1), CODE(0) => ALUCODE(0), 
                           DATA1(31) => MUXNPCout_31_port, DATA1(30) => 
                           MUXNPCout_30_port, DATA1(29) => MUXNPCout_29_port, 
                           DATA1(28) => MUXNPCout_28_port, DATA1(27) => 
                           MUXNPCout_27_port, DATA1(26) => MUXNPCout_26_port, 
                           DATA1(25) => MUXNPCout_25_port, DATA1(24) => 
                           MUXNPCout_24_port, DATA1(23) => MUXNPCout_23_port, 
                           DATA1(22) => MUXNPCout_22_port, DATA1(21) => 
                           MUXNPCout_21_port, DATA1(20) => MUXNPCout_20_port, 
                           DATA1(19) => MUXNPCout_19_port, DATA1(18) => 
                           MUXNPCout_18_port, DATA1(17) => MUXNPCout_17_port, 
                           DATA1(16) => MUXNPCout_16_port, DATA1(15) => 
                           MUXNPCout_15_port, DATA1(14) => MUXNPCout_14_port, 
                           DATA1(13) => MUXNPCout_13_port, DATA1(12) => 
                           MUXNPCout_12_port, DATA1(11) => MUXNPCout_11_port, 
                           DATA1(10) => MUXNPCout_10_port, DATA1(9) => 
                           MUXNPCout_9_port, DATA1(8) => MUXNPCout_8_port, 
                           DATA1(7) => MUXNPCout_7_port, DATA1(6) => 
                           MUXNPCout_6_port, DATA1(5) => MUXNPCout_5_port, 
                           DATA1(4) => MUXNPCout_4_port, DATA1(3) => 
                           MUXNPCout_3_port, DATA1(2) => MUXNPCout_2_port, 
                           DATA1(1) => MUXNPCout_1_port, DATA1(0) => 
                           MUXNPCout_0_port, DATA2(31) => MUXWITH4out_31_port, 
                           DATA2(30) => MUXWITH4out_30_port, DATA2(29) => 
                           MUXWITH4out_29_port, DATA2(28) => 
                           MUXWITH4out_28_port, DATA2(27) => 
                           MUXWITH4out_27_port, DATA2(26) => 
                           MUXWITH4out_26_port, DATA2(25) => 
                           MUXWITH4out_25_port, DATA2(24) => 
                           MUXWITH4out_24_port, DATA2(23) => 
                           MUXWITH4out_23_port, DATA2(22) => 
                           MUXWITH4out_22_port, DATA2(21) => 
                           MUXWITH4out_21_port, DATA2(20) => 
                           MUXWITH4out_20_port, DATA2(19) => 
                           MUXWITH4out_19_port, DATA2(18) => 
                           MUXWITH4out_18_port, DATA2(17) => 
                           MUXWITH4out_17_port, DATA2(16) => 
                           MUXWITH4out_16_port, DATA2(15) => 
                           MUXWITH4out_15_port, DATA2(14) => 
                           MUXWITH4out_14_port, DATA2(13) => 
                           MUXWITH4out_13_port, DATA2(12) => 
                           MUXWITH4out_12_port, DATA2(11) => 
                           MUXWITH4out_11_port, DATA2(10) => 
                           MUXWITH4out_10_port, DATA2(9) => MUXWITH4out_9_port,
                           DATA2(8) => MUXWITH4out_8_port, DATA2(7) => 
                           MUXWITH4out_7_port, DATA2(6) => MUXWITH4out_6_port, 
                           DATA2(5) => MUXWITH4out_5_port, DATA2(4) => 
                           MUXWITH4out_4_port, DATA2(3) => MUXWITH4out_3_port, 
                           DATA2(2) => MUXWITH4out_2_port, DATA2(1) => 
                           MUXWITH4out_1_port, DATA2(0) => MUXWITH4out_0_port, 
                           OUTALU(31) => ALUout_31_port, OUTALU(30) => 
                           ALUout_30_port, OUTALU(29) => ALUout_29_port, 
                           OUTALU(28) => ALUout_28_port, OUTALU(27) => 
                           ALUout_27_port, OUTALU(26) => ALUout_26_port, 
                           OUTALU(25) => ALUout_25_port, OUTALU(24) => 
                           ALUout_24_port, OUTALU(23) => ALUout_23_port, 
                           OUTALU(22) => ALUout_22_port, OUTALU(21) => 
                           ALUout_21_port, OUTALU(20) => ALUout_20_port, 
                           OUTALU(19) => ALUout_19_port, OUTALU(18) => 
                           ALUout_18_port, OUTALU(17) => ALUout_17_port, 
                           OUTALU(16) => ALUout_16_port, OUTALU(15) => 
                           ALUout_15_port, OUTALU(14) => ALUout_14_port, 
                           OUTALU(13) => ALUout_13_port, OUTALU(12) => 
                           ALUout_12_port, OUTALU(11) => ALUout_11_port, 
                           OUTALU(10) => ALUout_10_port, OUTALU(9) => 
                           ALUout_9_port, OUTALU(8) => ALUout_8_port, OUTALU(7)
                           => ALUout_7_port, OUTALU(6) => ALUout_6_port, 
                           OUTALU(5) => ALUout_5_port, OUTALU(4) => 
                           ALUout_4_port, OUTALU(3) => ALUout_3_port, OUTALU(2)
                           => ALUout_2_port, OUTALU(1) => ALUout_1_port, 
                           OUTALU(0) => ALUout_0_port);
   ALUout_REG : reg_6 port map( clock => clock, reset => reset, load => en3, 
                           i(31) => ALUout_31_port, i(30) => ALUout_30_port, 
                           i(29) => ALUout_29_port, i(28) => ALUout_28_port, 
                           i(27) => ALUout_27_port, i(26) => ALUout_26_port, 
                           i(25) => ALUout_25_port, i(24) => ALUout_24_port, 
                           i(23) => ALUout_23_port, i(22) => ALUout_22_port, 
                           i(21) => ALUout_21_port, i(20) => ALUout_20_port, 
                           i(19) => ALUout_19_port, i(18) => ALUout_18_port, 
                           i(17) => ALUout_17_port, i(16) => ALUout_16_port, 
                           i(15) => ALUout_15_port, i(14) => ALUout_14_port, 
                           i(13) => ALUout_13_port, i(12) => ALUout_12_port, 
                           i(11) => ALUout_11_port, i(10) => ALUout_10_port, 
                           i(9) => ALUout_9_port, i(8) => ALUout_8_port, i(7) 
                           => ALUout_7_port, i(6) => ALUout_6_port, i(5) => 
                           ALUout_5_port, i(4) => ALUout_4_port, i(3) => 
                           ALUout_3_port, i(2) => ALUout_2_port, i(1) => 
                           ALUout_1_port, i(0) => ALUout_0_port, o(31) => 
                           ALUtoMEMORY(31), o(30) => ALUtoMEMORY(30), o(29) => 
                           ALUtoMEMORY(29), o(28) => ALUtoMEMORY(28), o(27) => 
                           ALUtoMEMORY(27), o(26) => ALUtoMEMORY(26), o(25) => 
                           ALUtoMEMORY(25), o(24) => ALUtoMEMORY(24), o(23) => 
                           ALUtoMEMORY(23), o(22) => ALUtoMEMORY(22), o(21) => 
                           ALUtoMEMORY(21), o(20) => ALUtoMEMORY(20), o(19) => 
                           ALUtoMEMORY(19), o(18) => ALUtoMEMORY(18), o(17) => 
                           ALUtoMEMORY(17), o(16) => ALUtoMEMORY(16), o(15) => 
                           ALUtoMEMORY(15), o(14) => ALUtoMEMORY(14), o(13) => 
                           ALUtoMEMORY(13), o(12) => ALUtoMEMORY(12), o(11) => 
                           ALUtoMEMORY(11), o(10) => ALUtoMEMORY(10), o(9) => 
                           ALUtoMEMORY(9), o(8) => ALUtoMEMORY(8), o(7) => 
                           ALUtoMEMORY(7), o(6) => ALUtoMEMORY(6), o(5) => 
                           ALUtoMEMORY(5), o(4) => ALUtoMEMORY(4), o(3) => 
                           ALUtoMEMORY(3), o(2) => ALUtoMEMORY(2), o(1) => 
                           ALUtoMEMORY(1), o(0) => ALUtoMEMORY(0));
   RFout2_REG : reg_5 port map( clock => clock, reset => reset, load => en3, 
                           i(31) => OUT2RF(31), i(30) => OUT2RF(30), i(29) => 
                           OUT2RF(29), i(28) => OUT2RF(28), i(27) => OUT2RF(27)
                           , i(26) => OUT2RF(26), i(25) => OUT2RF(25), i(24) =>
                           OUT2RF(24), i(23) => OUT2RF(23), i(22) => OUT2RF(22)
                           , i(21) => OUT2RF(21), i(20) => OUT2RF(20), i(19) =>
                           OUT2RF(19), i(18) => OUT2RF(18), i(17) => OUT2RF(17)
                           , i(16) => OUT2RF(16), i(15) => OUT2RF(15), i(14) =>
                           OUT2RF(14), i(13) => OUT2RF(13), i(12) => OUT2RF(12)
                           , i(11) => OUT2RF(11), i(10) => OUT2RF(10), i(9) => 
                           OUT2RF(9), i(8) => OUT2RF(8), i(7) => OUT2RF(7), 
                           i(6) => OUT2RF(6), i(5) => OUT2RF(5), i(4) => 
                           OUT2RF(4), i(3) => OUT2RF(3), i(2) => OUT2RF(2), 
                           i(1) => OUT2RF(1), i(0) => OUT2RF(0), o(31) => 
                           OUT2RFtoMEMORY(31), o(30) => OUT2RFtoMEMORY(30), 
                           o(29) => OUT2RFtoMEMORY(29), o(28) => 
                           OUT2RFtoMEMORY(28), o(27) => OUT2RFtoMEMORY(27), 
                           o(26) => OUT2RFtoMEMORY(26), o(25) => 
                           OUT2RFtoMEMORY(25), o(24) => OUT2RFtoMEMORY(24), 
                           o(23) => OUT2RFtoMEMORY(23), o(22) => 
                           OUT2RFtoMEMORY(22), o(21) => OUT2RFtoMEMORY(21), 
                           o(20) => OUT2RFtoMEMORY(20), o(19) => 
                           OUT2RFtoMEMORY(19), o(18) => OUT2RFtoMEMORY(18), 
                           o(17) => OUT2RFtoMEMORY(17), o(16) => 
                           OUT2RFtoMEMORY(16), o(15) => OUT2RFtoMEMORY(15), 
                           o(14) => OUT2RFtoMEMORY(14), o(13) => 
                           OUT2RFtoMEMORY(13), o(12) => OUT2RFtoMEMORY(12), 
                           o(11) => OUT2RFtoMEMORY(11), o(10) => 
                           OUT2RFtoMEMORY(10), o(9) => OUT2RFtoMEMORY(9), o(8) 
                           => OUT2RFtoMEMORY(8), o(7) => OUT2RFtoMEMORY(7), 
                           o(6) => OUT2RFtoMEMORY(6), o(5) => OUT2RFtoMEMORY(5)
                           , o(4) => OUT2RFtoMEMORY(4), o(3) => 
                           OUT2RFtoMEMORY(3), o(2) => OUT2RFtoMEMORY(2), o(1) 
                           => OUT2RFtoMEMORY(1), o(0) => OUT2RFtoMEMORY(0));
   AddressW_REG : reg_4 port map( clock => clock, reset => reset, load => en3, 
                           i(31) => AddressWfromDecode(31), i(30) => 
                           AddressWfromDecode(30), i(29) => 
                           AddressWfromDecode(29), i(28) => 
                           AddressWfromDecode(28), i(27) => 
                           AddressWfromDecode(27), i(26) => 
                           AddressWfromDecode(26), i(25) => 
                           AddressWfromDecode(25), i(24) => 
                           AddressWfromDecode(24), i(23) => 
                           AddressWfromDecode(23), i(22) => 
                           AddressWfromDecode(22), i(21) => 
                           AddressWfromDecode(21), i(20) => 
                           AddressWfromDecode(20), i(19) => 
                           AddressWfromDecode(19), i(18) => 
                           AddressWfromDecode(18), i(17) => 
                           AddressWfromDecode(17), i(16) => 
                           AddressWfromDecode(16), i(15) => 
                           AddressWfromDecode(15), i(14) => 
                           AddressWfromDecode(14), i(13) => 
                           AddressWfromDecode(13), i(12) => 
                           AddressWfromDecode(12), i(11) => 
                           AddressWfromDecode(11), i(10) => 
                           AddressWfromDecode(10), i(9) => 
                           AddressWfromDecode(9), i(8) => AddressWfromDecode(8)
                           , i(7) => AddressWfromDecode(7), i(6) => 
                           AddressWfromDecode(6), i(5) => AddressWfromDecode(5)
                           , i(4) => AddressWfromDecode(4), i(3) => 
                           AddressWfromDecode(3), i(2) => AddressWfromDecode(2)
                           , i(1) => AddressWfromDecode(1), i(0) => 
                           AddressWfromDecode(0), o(31) => AddressWtoMEMORY(31)
                           , o(30) => AddressWtoMEMORY(30), o(29) => 
                           AddressWtoMEMORY(29), o(28) => AddressWtoMEMORY(28),
                           o(27) => AddressWtoMEMORY(27), o(26) => 
                           AddressWtoMEMORY(26), o(25) => AddressWtoMEMORY(25),
                           o(24) => AddressWtoMEMORY(24), o(23) => 
                           AddressWtoMEMORY(23), o(22) => AddressWtoMEMORY(22),
                           o(21) => AddressWtoMEMORY(21), o(20) => 
                           AddressWtoMEMORY(20), o(19) => AddressWtoMEMORY(19),
                           o(18) => AddressWtoMEMORY(18), o(17) => 
                           AddressWtoMEMORY(17), o(16) => AddressWtoMEMORY(16),
                           o(15) => AddressWtoMEMORY(15), o(14) => 
                           AddressWtoMEMORY(14), o(13) => AddressWtoMEMORY(13),
                           o(12) => AddressWtoMEMORY(12), o(11) => 
                           AddressWtoMEMORY(11), o(10) => AddressWtoMEMORY(10),
                           o(9) => AddressWtoMEMORY(9), o(8) => 
                           AddressWtoMEMORY(8), o(7) => AddressWtoMEMORY(7), 
                           o(6) => AddressWtoMEMORY(6), o(5) => 
                           AddressWtoMEMORY(5), o(4) => AddressWtoMEMORY(4), 
                           o(3) => AddressWtoMEMORY(3), o(2) => 
                           AddressWtoMEMORY(2), o(1) => AddressWtoMEMORY(1), 
                           o(0) => AddressWtoMEMORY(0));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity DecodeUnit is

   port( clock, reset, JMP, RegDestination, en2, SignSelect, BranchCondSel, 
         BRANCHenable, RD1, RD2, WR : in std_logic;  Instruction : in 
         std_logic_vector (31 downto 0);  ADD_WR : in std_logic_vector (4 
         downto 0);  DATAIN, NPCfromIF : in std_logic_vector (31 downto 0);  
         OUT1, OUT2, OUTNPC, OUTIMM, NPCtoEX, AddressWtoEX : out 
         std_logic_vector (31 downto 0);  BRANCHtoFetch : out std_logic);

end DecodeUnit;

architecture SYN_structural of DecodeUnit is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DecodeUnit_DW01_add_0
      port( A, B : in std_logic_vector (9 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (9 downto 0);  CO : out std_logic);
   end component;
   
   component register_file
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component reg_7
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_8
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_9
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_10
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_11
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component BranchUnit
      port( a : in std_logic_vector (31 downto 0);  sel : in std_logic;  y : 
            out std_logic);
   end component;
   
   component Mux21_5
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component Mux41
      port( a, b, c, d : in std_logic_vector (31 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  y : out std_logic_vector (31 downto
            0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, OUTNPC_9_port, OUTNPC_8_port, 
      OUTNPC_7_port, OUTNPC_6_port, OUTNPC_5_port, OUTNPC_4_port, OUTNPC_3_port
      , OUTNPC_2_port, OUTNPC_1_port, OUTNPC_0_port, AddressW_31_port, 
      AddressW_30_port, AddressW_29_port, AddressW_28_port, AddressW_27_port, 
      AddressW_26_port, AddressW_25_port, AddressW_24_port, AddressW_23_port, 
      AddressW_22_port, AddressW_21_port, AddressW_20_port, AddressW_19_port, 
      AddressW_18_port, AddressW_17_port, AddressW_16_port, AddressW_15_port, 
      AddressW_14_port, AddressW_13_port, AddressW_12_port, AddressW_11_port, 
      AddressW_10_port, AddressW_9_port, AddressW_8_port, AddressW_7_port, 
      AddressW_6_port, AddressW_5_port, AddressW_4_port, AddressW_3_port, 
      AddressW_2_port, AddressW_1_port, AddressW_0_port, MuxtoIMM_31_port, 
      MuxtoIMM_30_port, MuxtoIMM_29_port, MuxtoIMM_28_port, MuxtoIMM_27_port, 
      MuxtoIMM_26_port, MuxtoIMM_25_port, MuxtoIMM_24_port, MuxtoIMM_23_port, 
      MuxtoIMM_22_port, MuxtoIMM_21_port, MuxtoIMM_20_port, MuxtoIMM_19_port, 
      MuxtoIMM_18_port, MuxtoIMM_17_port, MuxtoIMM_16_port, MuxtoIMM_15_port, 
      MuxtoIMM_14_port, MuxtoIMM_13_port, MuxtoIMM_12_port, MuxtoIMM_11_port, 
      MuxtoIMM_10_port, MuxtoIMM_9_port, MuxtoIMM_8_port, MuxtoIMM_7_port, 
      MuxtoIMM_6_port, MuxtoIMM_5_port, MuxtoIMM_4_port, MuxtoIMM_3_port, 
      MuxtoIMM_2_port, MuxtoIMM_1_port, MuxtoIMM_0_port, RFOUT1_31_port, 
      RFOUT1_30_port, RFOUT1_29_port, RFOUT1_28_port, RFOUT1_27_port, 
      RFOUT1_26_port, RFOUT1_25_port, RFOUT1_24_port, RFOUT1_23_port, 
      RFOUT1_22_port, RFOUT1_21_port, RFOUT1_20_port, RFOUT1_19_port, 
      RFOUT1_18_port, RFOUT1_17_port, RFOUT1_16_port, RFOUT1_15_port, 
      RFOUT1_14_port, RFOUT1_13_port, RFOUT1_12_port, RFOUT1_11_port, 
      RFOUT1_10_port, RFOUT1_9_port, RFOUT1_8_port, RFOUT1_7_port, 
      RFOUT1_6_port, RFOUT1_5_port, RFOUT1_4_port, RFOUT1_3_port, RFOUT1_2_port
      , RFOUT1_1_port, RFOUT1_0_port, BranchTaken, RFOUT2_31_port, 
      RFOUT2_30_port, RFOUT2_29_port, RFOUT2_28_port, RFOUT2_27_port, 
      RFOUT2_26_port, RFOUT2_25_port, RFOUT2_24_port, RFOUT2_23_port, 
      RFOUT2_22_port, RFOUT2_21_port, RFOUT2_20_port, RFOUT2_19_port, 
      RFOUT2_18_port, RFOUT2_17_port, RFOUT2_16_port, RFOUT2_15_port, 
      RFOUT2_14_port, RFOUT2_13_port, RFOUT2_12_port, RFOUT2_11_port, 
      RFOUT2_10_port, RFOUT2_9_port, RFOUT2_8_port, RFOUT2_7_port, 
      RFOUT2_6_port, RFOUT2_5_port, RFOUT2_4_port, RFOUT2_3_port, RFOUT2_2_port
      , RFOUT2_1_port, RFOUT2_0_port, n2, n4, n20, n_1352 : std_logic;

begin
   OUTNPC <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port
      , X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      OUTNPC_9_port, OUTNPC_8_port, OUTNPC_7_port, OUTNPC_6_port, OUTNPC_5_port
      , OUTNPC_4_port, OUTNPC_3_port, OUTNPC_2_port, OUTNPC_1_port, 
      OUTNPC_0_port );
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n2 <= '0';
   ADDRESS_MUX : Mux41 port map( a(31) => X_Logic0_port, a(30) => X_Logic0_port
                           , a(29) => X_Logic0_port, a(28) => X_Logic0_port, 
                           a(27) => X_Logic0_port, a(26) => X_Logic0_port, 
                           a(25) => X_Logic0_port, a(24) => X_Logic0_port, 
                           a(23) => X_Logic0_port, a(22) => X_Logic0_port, 
                           a(21) => X_Logic0_port, a(20) => X_Logic0_port, 
                           a(19) => X_Logic0_port, a(18) => X_Logic0_port, 
                           a(17) => X_Logic0_port, a(16) => X_Logic0_port, 
                           a(15) => X_Logic0_port, a(14) => X_Logic0_port, 
                           a(13) => X_Logic0_port, a(12) => X_Logic0_port, 
                           a(11) => X_Logic0_port, a(10) => X_Logic0_port, a(9)
                           => X_Logic0_port, a(8) => X_Logic0_port, a(7) => 
                           X_Logic0_port, a(6) => X_Logic0_port, a(5) => 
                           X_Logic0_port, a(4) => Instruction(20), a(3) => 
                           Instruction(19), a(2) => Instruction(18), a(1) => 
                           Instruction(17), a(0) => Instruction(16), b(31) => 
                           X_Logic0_port, b(30) => X_Logic0_port, b(29) => 
                           X_Logic0_port, b(28) => X_Logic0_port, b(27) => 
                           X_Logic0_port, b(26) => X_Logic0_port, b(25) => 
                           X_Logic0_port, b(24) => X_Logic0_port, b(23) => 
                           X_Logic0_port, b(22) => X_Logic0_port, b(21) => 
                           X_Logic0_port, b(20) => X_Logic0_port, b(19) => 
                           X_Logic0_port, b(18) => X_Logic0_port, b(17) => 
                           X_Logic0_port, b(16) => X_Logic0_port, b(15) => 
                           X_Logic0_port, b(14) => X_Logic0_port, b(13) => 
                           X_Logic0_port, b(12) => X_Logic0_port, b(11) => 
                           X_Logic0_port, b(10) => X_Logic0_port, b(9) => 
                           X_Logic0_port, b(8) => X_Logic0_port, b(7) => 
                           X_Logic0_port, b(6) => X_Logic0_port, b(5) => 
                           X_Logic0_port, b(4) => Instruction(15), b(3) => 
                           Instruction(14), b(2) => Instruction(13), b(1) => 
                           Instruction(12), b(0) => Instruction(11), c(31) => 
                           X_Logic0_port, c(30) => X_Logic0_port, c(29) => 
                           X_Logic0_port, c(28) => X_Logic0_port, c(27) => 
                           X_Logic0_port, c(26) => X_Logic0_port, c(25) => 
                           X_Logic0_port, c(24) => X_Logic0_port, c(23) => 
                           X_Logic0_port, c(22) => X_Logic0_port, c(21) => 
                           X_Logic0_port, c(20) => X_Logic0_port, c(19) => 
                           X_Logic0_port, c(18) => X_Logic0_port, c(17) => 
                           X_Logic0_port, c(16) => X_Logic0_port, c(15) => 
                           X_Logic0_port, c(14) => X_Logic0_port, c(13) => 
                           X_Logic0_port, c(12) => X_Logic0_port, c(11) => 
                           X_Logic0_port, c(10) => X_Logic0_port, c(9) => 
                           X_Logic0_port, c(8) => X_Logic0_port, c(7) => 
                           X_Logic0_port, c(6) => X_Logic0_port, c(5) => 
                           X_Logic0_port, c(4) => X_Logic1_port, c(3) => 
                           X_Logic1_port, c(2) => X_Logic1_port, c(1) => 
                           X_Logic1_port, c(0) => X_Logic1_port, d(31) => 
                           X_Logic0_port, d(30) => X_Logic0_port, d(29) => 
                           X_Logic0_port, d(28) => X_Logic0_port, d(27) => 
                           X_Logic0_port, d(26) => X_Logic0_port, d(25) => 
                           X_Logic0_port, d(24) => X_Logic0_port, d(23) => 
                           X_Logic0_port, d(22) => X_Logic0_port, d(21) => 
                           X_Logic0_port, d(20) => X_Logic0_port, d(19) => 
                           X_Logic0_port, d(18) => X_Logic0_port, d(17) => 
                           X_Logic0_port, d(16) => X_Logic0_port, d(15) => 
                           X_Logic0_port, d(14) => X_Logic0_port, d(13) => 
                           X_Logic0_port, d(12) => X_Logic0_port, d(11) => 
                           X_Logic0_port, d(10) => X_Logic0_port, d(9) => 
                           X_Logic0_port, d(8) => X_Logic0_port, d(7) => 
                           X_Logic0_port, d(6) => X_Logic0_port, d(5) => 
                           X_Logic0_port, d(4) => X_Logic1_port, d(3) => 
                           X_Logic1_port, d(2) => X_Logic1_port, d(1) => 
                           X_Logic1_port, d(0) => X_Logic1_port, sel(1) => JMP,
                           sel(0) => RegDestination, y(31) => AddressW_31_port,
                           y(30) => AddressW_30_port, y(29) => AddressW_29_port
                           , y(28) => AddressW_28_port, y(27) => 
                           AddressW_27_port, y(26) => AddressW_26_port, y(25) 
                           => AddressW_25_port, y(24) => AddressW_24_port, 
                           y(23) => AddressW_23_port, y(22) => AddressW_22_port
                           , y(21) => AddressW_21_port, y(20) => 
                           AddressW_20_port, y(19) => AddressW_19_port, y(18) 
                           => AddressW_18_port, y(17) => AddressW_17_port, 
                           y(16) => AddressW_16_port, y(15) => AddressW_15_port
                           , y(14) => AddressW_14_port, y(13) => 
                           AddressW_13_port, y(12) => AddressW_12_port, y(11) 
                           => AddressW_11_port, y(10) => AddressW_10_port, y(9)
                           => AddressW_9_port, y(8) => AddressW_8_port, y(7) =>
                           AddressW_7_port, y(6) => AddressW_6_port, y(5) => 
                           AddressW_5_port, y(4) => AddressW_4_port, y(3) => 
                           AddressW_3_port, y(2) => AddressW_2_port, y(1) => 
                           AddressW_1_port, y(0) => AddressW_0_port);
   MUX : Mux21_5 port map( a(31) => Instruction(15), a(30) => Instruction(15), 
                           a(29) => Instruction(15), a(28) => Instruction(15), 
                           a(27) => Instruction(15), a(26) => Instruction(15), 
                           a(25) => Instruction(15), a(24) => Instruction(15), 
                           a(23) => Instruction(15), a(22) => Instruction(15), 
                           a(21) => Instruction(15), a(20) => Instruction(15), 
                           a(19) => Instruction(15), a(18) => Instruction(15), 
                           a(17) => Instruction(15), a(16) => Instruction(15), 
                           a(15) => Instruction(15), a(14) => Instruction(14), 
                           a(13) => Instruction(13), a(12) => Instruction(12), 
                           a(11) => Instruction(11), a(10) => Instruction(10), 
                           a(9) => Instruction(9), a(8) => Instruction(8), a(7)
                           => Instruction(7), a(6) => Instruction(6), a(5) => 
                           Instruction(5), a(4) => Instruction(4), a(3) => 
                           Instruction(3), a(2) => Instruction(2), a(1) => 
                           Instruction(1), a(0) => Instruction(0), b(31) => n20
                           , b(30) => n20, b(29) => n20, b(28) => n20, b(27) =>
                           n20, b(26) => n20, b(25) => n20, b(24) => 
                           Instruction(24), b(23) => Instruction(23), b(22) => 
                           Instruction(22), b(21) => Instruction(21), b(20) => 
                           Instruction(20), b(19) => Instruction(19), b(18) => 
                           Instruction(18), b(17) => Instruction(17), b(16) => 
                           Instruction(16), b(15) => Instruction(15), b(14) => 
                           Instruction(14), b(13) => Instruction(13), b(12) => 
                           Instruction(12), b(11) => Instruction(11), b(10) => 
                           Instruction(10), b(9) => Instruction(9), b(8) => 
                           Instruction(8), b(7) => Instruction(7), b(6) => 
                           Instruction(6), b(5) => Instruction(5), b(4) => 
                           Instruction(4), b(3) => Instruction(3), b(2) => 
                           Instruction(2), b(1) => Instruction(1), b(0) => 
                           Instruction(0), sel => SignSelect, y(31) => 
                           MuxtoIMM_31_port, y(30) => MuxtoIMM_30_port, y(29) 
                           => MuxtoIMM_29_port, y(28) => MuxtoIMM_28_port, 
                           y(27) => MuxtoIMM_27_port, y(26) => MuxtoIMM_26_port
                           , y(25) => MuxtoIMM_25_port, y(24) => 
                           MuxtoIMM_24_port, y(23) => MuxtoIMM_23_port, y(22) 
                           => MuxtoIMM_22_port, y(21) => MuxtoIMM_21_port, 
                           y(20) => MuxtoIMM_20_port, y(19) => MuxtoIMM_19_port
                           , y(18) => MuxtoIMM_18_port, y(17) => 
                           MuxtoIMM_17_port, y(16) => MuxtoIMM_16_port, y(15) 
                           => MuxtoIMM_15_port, y(14) => MuxtoIMM_14_port, 
                           y(13) => MuxtoIMM_13_port, y(12) => MuxtoIMM_12_port
                           , y(11) => MuxtoIMM_11_port, y(10) => 
                           MuxtoIMM_10_port, y(9) => MuxtoIMM_9_port, y(8) => 
                           MuxtoIMM_8_port, y(7) => MuxtoIMM_7_port, y(6) => 
                           MuxtoIMM_6_port, y(5) => MuxtoIMM_5_port, y(4) => 
                           MuxtoIMM_4_port, y(3) => MuxtoIMM_3_port, y(2) => 
                           MuxtoIMM_2_port, y(1) => MuxtoIMM_1_port, y(0) => 
                           MuxtoIMM_0_port);
   BRANCH : BranchUnit port map( a(31) => RFOUT1_31_port, a(30) => 
                           RFOUT1_30_port, a(29) => RFOUT1_29_port, a(28) => 
                           RFOUT1_28_port, a(27) => RFOUT1_27_port, a(26) => 
                           RFOUT1_26_port, a(25) => RFOUT1_25_port, a(24) => 
                           RFOUT1_24_port, a(23) => RFOUT1_23_port, a(22) => 
                           RFOUT1_22_port, a(21) => RFOUT1_21_port, a(20) => 
                           RFOUT1_20_port, a(19) => RFOUT1_19_port, a(18) => 
                           RFOUT1_18_port, a(17) => RFOUT1_17_port, a(16) => 
                           RFOUT1_16_port, a(15) => RFOUT1_15_port, a(14) => 
                           RFOUT1_14_port, a(13) => RFOUT1_13_port, a(12) => 
                           RFOUT1_12_port, a(11) => RFOUT1_11_port, a(10) => 
                           RFOUT1_10_port, a(9) => RFOUT1_9_port, a(8) => 
                           RFOUT1_8_port, a(7) => RFOUT1_7_port, a(6) => 
                           RFOUT1_6_port, a(5) => RFOUT1_5_port, a(4) => 
                           RFOUT1_4_port, a(3) => RFOUT1_3_port, a(2) => 
                           RFOUT1_2_port, a(1) => RFOUT1_1_port, a(0) => 
                           RFOUT1_0_port, sel => BranchCondSel, y => 
                           BranchTaken);
   IMM_REG : reg_11 port map( clock => clock, reset => reset, load => en2, 
                           i(31) => MuxtoIMM_31_port, i(30) => MuxtoIMM_30_port
                           , i(29) => MuxtoIMM_29_port, i(28) => 
                           MuxtoIMM_28_port, i(27) => MuxtoIMM_27_port, i(26) 
                           => MuxtoIMM_26_port, i(25) => MuxtoIMM_25_port, 
                           i(24) => MuxtoIMM_24_port, i(23) => MuxtoIMM_23_port
                           , i(22) => MuxtoIMM_22_port, i(21) => 
                           MuxtoIMM_21_port, i(20) => MuxtoIMM_20_port, i(19) 
                           => MuxtoIMM_19_port, i(18) => MuxtoIMM_18_port, 
                           i(17) => MuxtoIMM_17_port, i(16) => MuxtoIMM_16_port
                           , i(15) => MuxtoIMM_15_port, i(14) => 
                           MuxtoIMM_14_port, i(13) => MuxtoIMM_13_port, i(12) 
                           => MuxtoIMM_12_port, i(11) => MuxtoIMM_11_port, 
                           i(10) => MuxtoIMM_10_port, i(9) => MuxtoIMM_9_port, 
                           i(8) => MuxtoIMM_8_port, i(7) => MuxtoIMM_7_port, 
                           i(6) => MuxtoIMM_6_port, i(5) => MuxtoIMM_5_port, 
                           i(4) => MuxtoIMM_4_port, i(3) => MuxtoIMM_3_port, 
                           i(2) => MuxtoIMM_2_port, i(1) => MuxtoIMM_1_port, 
                           i(0) => MuxtoIMM_0_port, o(31) => OUTIMM(31), o(30) 
                           => OUTIMM(30), o(29) => OUTIMM(29), o(28) => 
                           OUTIMM(28), o(27) => OUTIMM(27), o(26) => OUTIMM(26)
                           , o(25) => OUTIMM(25), o(24) => OUTIMM(24), o(23) =>
                           OUTIMM(23), o(22) => OUTIMM(22), o(21) => OUTIMM(21)
                           , o(20) => OUTIMM(20), o(19) => OUTIMM(19), o(18) =>
                           OUTIMM(18), o(17) => OUTIMM(17), o(16) => OUTIMM(16)
                           , o(15) => OUTIMM(15), o(14) => OUTIMM(14), o(13) =>
                           OUTIMM(13), o(12) => OUTIMM(12), o(11) => OUTIMM(11)
                           , o(10) => OUTIMM(10), o(9) => OUTIMM(9), o(8) => 
                           OUTIMM(8), o(7) => OUTIMM(7), o(6) => OUTIMM(6), 
                           o(5) => OUTIMM(5), o(4) => OUTIMM(4), o(3) => 
                           OUTIMM(3), o(2) => OUTIMM(2), o(1) => OUTIMM(1), 
                           o(0) => OUTIMM(0));
   OUT1_REG : reg_10 port map( clock => clock, reset => reset, load => en2, 
                           i(31) => RFOUT1_31_port, i(30) => RFOUT1_30_port, 
                           i(29) => RFOUT1_29_port, i(28) => RFOUT1_28_port, 
                           i(27) => RFOUT1_27_port, i(26) => RFOUT1_26_port, 
                           i(25) => RFOUT1_25_port, i(24) => RFOUT1_24_port, 
                           i(23) => RFOUT1_23_port, i(22) => RFOUT1_22_port, 
                           i(21) => RFOUT1_21_port, i(20) => RFOUT1_20_port, 
                           i(19) => RFOUT1_19_port, i(18) => RFOUT1_18_port, 
                           i(17) => RFOUT1_17_port, i(16) => RFOUT1_16_port, 
                           i(15) => RFOUT1_15_port, i(14) => RFOUT1_14_port, 
                           i(13) => RFOUT1_13_port, i(12) => RFOUT1_12_port, 
                           i(11) => RFOUT1_11_port, i(10) => RFOUT1_10_port, 
                           i(9) => RFOUT1_9_port, i(8) => RFOUT1_8_port, i(7) 
                           => RFOUT1_7_port, i(6) => RFOUT1_6_port, i(5) => 
                           RFOUT1_5_port, i(4) => RFOUT1_4_port, i(3) => 
                           RFOUT1_3_port, i(2) => RFOUT1_2_port, i(1) => 
                           RFOUT1_1_port, i(0) => RFOUT1_0_port, o(31) => 
                           OUT1(31), o(30) => OUT1(30), o(29) => OUT1(29), 
                           o(28) => OUT1(28), o(27) => OUT1(27), o(26) => 
                           OUT1(26), o(25) => OUT1(25), o(24) => OUT1(24), 
                           o(23) => OUT1(23), o(22) => OUT1(22), o(21) => 
                           OUT1(21), o(20) => OUT1(20), o(19) => OUT1(19), 
                           o(18) => OUT1(18), o(17) => OUT1(17), o(16) => 
                           OUT1(16), o(15) => OUT1(15), o(14) => OUT1(14), 
                           o(13) => OUT1(13), o(12) => OUT1(12), o(11) => 
                           OUT1(11), o(10) => OUT1(10), o(9) => OUT1(9), o(8) 
                           => OUT1(8), o(7) => OUT1(7), o(6) => OUT1(6), o(5) 
                           => OUT1(5), o(4) => OUT1(4), o(3) => OUT1(3), o(2) 
                           => OUT1(2), o(1) => OUT1(1), o(0) => OUT1(0));
   OUT2_REG : reg_9 port map( clock => clock, reset => reset, load => en2, 
                           i(31) => RFOUT2_31_port, i(30) => RFOUT2_30_port, 
                           i(29) => RFOUT2_29_port, i(28) => RFOUT2_28_port, 
                           i(27) => RFOUT2_27_port, i(26) => RFOUT2_26_port, 
                           i(25) => RFOUT2_25_port, i(24) => RFOUT2_24_port, 
                           i(23) => RFOUT2_23_port, i(22) => RFOUT2_22_port, 
                           i(21) => RFOUT2_21_port, i(20) => RFOUT2_20_port, 
                           i(19) => RFOUT2_19_port, i(18) => RFOUT2_18_port, 
                           i(17) => RFOUT2_17_port, i(16) => RFOUT2_16_port, 
                           i(15) => RFOUT2_15_port, i(14) => RFOUT2_14_port, 
                           i(13) => RFOUT2_13_port, i(12) => RFOUT2_12_port, 
                           i(11) => RFOUT2_11_port, i(10) => RFOUT2_10_port, 
                           i(9) => RFOUT2_9_port, i(8) => RFOUT2_8_port, i(7) 
                           => RFOUT2_7_port, i(6) => RFOUT2_6_port, i(5) => 
                           RFOUT2_5_port, i(4) => RFOUT2_4_port, i(3) => 
                           RFOUT2_3_port, i(2) => RFOUT2_2_port, i(1) => 
                           RFOUT2_1_port, i(0) => RFOUT2_0_port, o(31) => 
                           OUT2(31), o(30) => OUT2(30), o(29) => OUT2(29), 
                           o(28) => OUT2(28), o(27) => OUT2(27), o(26) => 
                           OUT2(26), o(25) => OUT2(25), o(24) => OUT2(24), 
                           o(23) => OUT2(23), o(22) => OUT2(22), o(21) => 
                           OUT2(21), o(20) => OUT2(20), o(19) => OUT2(19), 
                           o(18) => OUT2(18), o(17) => OUT2(17), o(16) => 
                           OUT2(16), o(15) => OUT2(15), o(14) => OUT2(14), 
                           o(13) => OUT2(13), o(12) => OUT2(12), o(11) => 
                           OUT2(11), o(10) => OUT2(10), o(9) => OUT2(9), o(8) 
                           => OUT2(8), o(7) => OUT2(7), o(6) => OUT2(6), o(5) 
                           => OUT2(5), o(4) => OUT2(4), o(3) => OUT2(3), o(2) 
                           => OUT2(2), o(1) => OUT2(1), o(0) => OUT2(0));
   NXPC_REG : reg_8 port map( clock => clock, reset => reset, load => en2, 
                           i(31) => NPCfromIF(31), i(30) => NPCfromIF(30), 
                           i(29) => NPCfromIF(29), i(28) => NPCfromIF(28), 
                           i(27) => NPCfromIF(27), i(26) => NPCfromIF(26), 
                           i(25) => NPCfromIF(25), i(24) => NPCfromIF(24), 
                           i(23) => NPCfromIF(23), i(22) => NPCfromIF(22), 
                           i(21) => NPCfromIF(21), i(20) => NPCfromIF(20), 
                           i(19) => NPCfromIF(19), i(18) => NPCfromIF(18), 
                           i(17) => NPCfromIF(17), i(16) => NPCfromIF(16), 
                           i(15) => NPCfromIF(15), i(14) => NPCfromIF(14), 
                           i(13) => NPCfromIF(13), i(12) => NPCfromIF(12), 
                           i(11) => NPCfromIF(11), i(10) => NPCfromIF(10), i(9)
                           => NPCfromIF(9), i(8) => NPCfromIF(8), i(7) => 
                           NPCfromIF(7), i(6) => NPCfromIF(6), i(5) => 
                           NPCfromIF(5), i(4) => NPCfromIF(4), i(3) => 
                           NPCfromIF(3), i(2) => NPCfromIF(2), i(1) => 
                           NPCfromIF(1), i(0) => NPCfromIF(0), o(31) => 
                           NPCtoEX(31), o(30) => NPCtoEX(30), o(29) => 
                           NPCtoEX(29), o(28) => NPCtoEX(28), o(27) => 
                           NPCtoEX(27), o(26) => NPCtoEX(26), o(25) => 
                           NPCtoEX(25), o(24) => NPCtoEX(24), o(23) => 
                           NPCtoEX(23), o(22) => NPCtoEX(22), o(21) => 
                           NPCtoEX(21), o(20) => NPCtoEX(20), o(19) => 
                           NPCtoEX(19), o(18) => NPCtoEX(18), o(17) => 
                           NPCtoEX(17), o(16) => NPCtoEX(16), o(15) => 
                           NPCtoEX(15), o(14) => NPCtoEX(14), o(13) => 
                           NPCtoEX(13), o(12) => NPCtoEX(12), o(11) => 
                           NPCtoEX(11), o(10) => NPCtoEX(10), o(9) => 
                           NPCtoEX(9), o(8) => NPCtoEX(8), o(7) => NPCtoEX(7), 
                           o(6) => NPCtoEX(6), o(5) => NPCtoEX(5), o(4) => 
                           NPCtoEX(4), o(3) => NPCtoEX(3), o(2) => NPCtoEX(2), 
                           o(1) => NPCtoEX(1), o(0) => NPCtoEX(0));
   ADD_WR_REG : reg_7 port map( clock => clock, reset => reset, load => en2, 
                           i(31) => AddressW_31_port, i(30) => AddressW_30_port
                           , i(29) => AddressW_29_port, i(28) => 
                           AddressW_28_port, i(27) => AddressW_27_port, i(26) 
                           => AddressW_26_port, i(25) => AddressW_25_port, 
                           i(24) => AddressW_24_port, i(23) => AddressW_23_port
                           , i(22) => AddressW_22_port, i(21) => 
                           AddressW_21_port, i(20) => AddressW_20_port, i(19) 
                           => AddressW_19_port, i(18) => AddressW_18_port, 
                           i(17) => AddressW_17_port, i(16) => AddressW_16_port
                           , i(15) => AddressW_15_port, i(14) => 
                           AddressW_14_port, i(13) => AddressW_13_port, i(12) 
                           => AddressW_12_port, i(11) => AddressW_11_port, 
                           i(10) => AddressW_10_port, i(9) => AddressW_9_port, 
                           i(8) => AddressW_8_port, i(7) => AddressW_7_port, 
                           i(6) => AddressW_6_port, i(5) => AddressW_5_port, 
                           i(4) => AddressW_4_port, i(3) => AddressW_3_port, 
                           i(2) => AddressW_2_port, i(1) => AddressW_1_port, 
                           i(0) => AddressW_0_port, o(31) => AddressWtoEX(31), 
                           o(30) => AddressWtoEX(30), o(29) => AddressWtoEX(29)
                           , o(28) => AddressWtoEX(28), o(27) => 
                           AddressWtoEX(27), o(26) => AddressWtoEX(26), o(25) 
                           => AddressWtoEX(25), o(24) => AddressWtoEX(24), 
                           o(23) => AddressWtoEX(23), o(22) => AddressWtoEX(22)
                           , o(21) => AddressWtoEX(21), o(20) => 
                           AddressWtoEX(20), o(19) => AddressWtoEX(19), o(18) 
                           => AddressWtoEX(18), o(17) => AddressWtoEX(17), 
                           o(16) => AddressWtoEX(16), o(15) => AddressWtoEX(15)
                           , o(14) => AddressWtoEX(14), o(13) => 
                           AddressWtoEX(13), o(12) => AddressWtoEX(12), o(11) 
                           => AddressWtoEX(11), o(10) => AddressWtoEX(10), o(9)
                           => AddressWtoEX(9), o(8) => AddressWtoEX(8), o(7) =>
                           AddressWtoEX(7), o(6) => AddressWtoEX(6), o(5) => 
                           AddressWtoEX(5), o(4) => AddressWtoEX(4), o(3) => 
                           AddressWtoEX(3), o(2) => AddressWtoEX(2), o(1) => 
                           AddressWtoEX(1), o(0) => AddressWtoEX(0));
   RF : register_file port map( CLK => clock, RESET => reset, ENABLE => 
                           X_Logic1_port, RD1 => RD1, RD2 => RD2, WR => WR, 
                           ADD_WR(4) => ADD_WR(4), ADD_WR(3) => ADD_WR(3), 
                           ADD_WR(2) => ADD_WR(2), ADD_WR(1) => ADD_WR(1), 
                           ADD_WR(0) => ADD_WR(0), ADD_RD1(4) => 
                           Instruction(25), ADD_RD1(3) => Instruction(24), 
                           ADD_RD1(2) => Instruction(23), ADD_RD1(1) => 
                           Instruction(22), ADD_RD1(0) => Instruction(21), 
                           ADD_RD2(4) => Instruction(20), ADD_RD2(3) => 
                           Instruction(19), ADD_RD2(2) => Instruction(18), 
                           ADD_RD2(1) => Instruction(17), ADD_RD2(0) => 
                           Instruction(16), DATAIN(31) => DATAIN(31), 
                           DATAIN(30) => DATAIN(30), DATAIN(29) => DATAIN(29), 
                           DATAIN(28) => DATAIN(28), DATAIN(27) => DATAIN(27), 
                           DATAIN(26) => DATAIN(26), DATAIN(25) => DATAIN(25), 
                           DATAIN(24) => DATAIN(24), DATAIN(23) => DATAIN(23), 
                           DATAIN(22) => DATAIN(22), DATAIN(21) => DATAIN(21), 
                           DATAIN(20) => DATAIN(20), DATAIN(19) => DATAIN(19), 
                           DATAIN(18) => DATAIN(18), DATAIN(17) => DATAIN(17), 
                           DATAIN(16) => DATAIN(16), DATAIN(15) => DATAIN(15), 
                           DATAIN(14) => DATAIN(14), DATAIN(13) => DATAIN(13), 
                           DATAIN(12) => DATAIN(12), DATAIN(11) => DATAIN(11), 
                           DATAIN(10) => DATAIN(10), DATAIN(9) => DATAIN(9), 
                           DATAIN(8) => DATAIN(8), DATAIN(7) => DATAIN(7), 
                           DATAIN(6) => DATAIN(6), DATAIN(5) => DATAIN(5), 
                           DATAIN(4) => DATAIN(4), DATAIN(3) => DATAIN(3), 
                           DATAIN(2) => DATAIN(2), DATAIN(1) => DATAIN(1), 
                           DATAIN(0) => DATAIN(0), OUT1(31) => RFOUT1_31_port, 
                           OUT1(30) => RFOUT1_30_port, OUT1(29) => 
                           RFOUT1_29_port, OUT1(28) => RFOUT1_28_port, OUT1(27)
                           => RFOUT1_27_port, OUT1(26) => RFOUT1_26_port, 
                           OUT1(25) => RFOUT1_25_port, OUT1(24) => 
                           RFOUT1_24_port, OUT1(23) => RFOUT1_23_port, OUT1(22)
                           => RFOUT1_22_port, OUT1(21) => RFOUT1_21_port, 
                           OUT1(20) => RFOUT1_20_port, OUT1(19) => 
                           RFOUT1_19_port, OUT1(18) => RFOUT1_18_port, OUT1(17)
                           => RFOUT1_17_port, OUT1(16) => RFOUT1_16_port, 
                           OUT1(15) => RFOUT1_15_port, OUT1(14) => 
                           RFOUT1_14_port, OUT1(13) => RFOUT1_13_port, OUT1(12)
                           => RFOUT1_12_port, OUT1(11) => RFOUT1_11_port, 
                           OUT1(10) => RFOUT1_10_port, OUT1(9) => RFOUT1_9_port
                           , OUT1(8) => RFOUT1_8_port, OUT1(7) => RFOUT1_7_port
                           , OUT1(6) => RFOUT1_6_port, OUT1(5) => RFOUT1_5_port
                           , OUT1(4) => RFOUT1_4_port, OUT1(3) => RFOUT1_3_port
                           , OUT1(2) => RFOUT1_2_port, OUT1(1) => RFOUT1_1_port
                           , OUT1(0) => RFOUT1_0_port, OUT2(31) => 
                           RFOUT2_31_port, OUT2(30) => RFOUT2_30_port, OUT2(29)
                           => RFOUT2_29_port, OUT2(28) => RFOUT2_28_port, 
                           OUT2(27) => RFOUT2_27_port, OUT2(26) => 
                           RFOUT2_26_port, OUT2(25) => RFOUT2_25_port, OUT2(24)
                           => RFOUT2_24_port, OUT2(23) => RFOUT2_23_port, 
                           OUT2(22) => RFOUT2_22_port, OUT2(21) => 
                           RFOUT2_21_port, OUT2(20) => RFOUT2_20_port, OUT2(19)
                           => RFOUT2_19_port, OUT2(18) => RFOUT2_18_port, 
                           OUT2(17) => RFOUT2_17_port, OUT2(16) => 
                           RFOUT2_16_port, OUT2(15) => RFOUT2_15_port, OUT2(14)
                           => RFOUT2_14_port, OUT2(13) => RFOUT2_13_port, 
                           OUT2(12) => RFOUT2_12_port, OUT2(11) => 
                           RFOUT2_11_port, OUT2(10) => RFOUT2_10_port, OUT2(9) 
                           => RFOUT2_9_port, OUT2(8) => RFOUT2_8_port, OUT2(7) 
                           => RFOUT2_7_port, OUT2(6) => RFOUT2_6_port, OUT2(5) 
                           => RFOUT2_5_port, OUT2(4) => RFOUT2_4_port, OUT2(3) 
                           => RFOUT2_3_port, OUT2(2) => RFOUT2_2_port, OUT2(1) 
                           => RFOUT2_1_port, OUT2(0) => RFOUT2_0_port);
   add_142 : DecodeUnit_DW01_add_0 port map( A(9) => NPCfromIF(9), A(8) => 
                           NPCfromIF(8), A(7) => NPCfromIF(7), A(6) => 
                           NPCfromIF(6), A(5) => NPCfromIF(5), A(4) => 
                           NPCfromIF(4), A(3) => NPCfromIF(3), A(2) => 
                           NPCfromIF(2), A(1) => NPCfromIF(1), A(0) => 
                           NPCfromIF(0), B(9) => MuxtoIMM_11_port, B(8) => 
                           MuxtoIMM_10_port, B(7) => MuxtoIMM_9_port, B(6) => 
                           MuxtoIMM_8_port, B(5) => MuxtoIMM_7_port, B(4) => 
                           MuxtoIMM_6_port, B(3) => MuxtoIMM_5_port, B(2) => 
                           MuxtoIMM_4_port, B(1) => MuxtoIMM_3_port, B(0) => 
                           MuxtoIMM_2_port, CI => n2, SUM(9) => OUTNPC_9_port, 
                           SUM(8) => OUTNPC_8_port, SUM(7) => OUTNPC_7_port, 
                           SUM(6) => OUTNPC_6_port, SUM(5) => OUTNPC_5_port, 
                           SUM(4) => OUTNPC_4_port, SUM(3) => OUTNPC_3_port, 
                           SUM(2) => OUTNPC_2_port, SUM(1) => OUTNPC_1_port, 
                           SUM(0) => OUTNPC_0_port, CO => n_1352);
   U3 : INV_X1 port map( A => n4, ZN => BRANCHtoFetch);
   U5 : CLKBUF_X1 port map( A => Instruction(25), Z => n20);
   U6 : AOI21_X1 port map( B1 => BranchTaken, B2 => BRANCHenable, A => JMP, ZN 
                           => n4);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity fetchUnit is

   port( clock, reset, en1 : in std_logic;  BranchPC : in std_logic_vector (31 
         downto 0);  BRANCHfromDECODE : in std_logic;  Instruction : in 
         std_logic_vector (31 downto 0);  PCtoIM, IRtoDecode, NPCtoDecode : out
         std_logic_vector (31 downto 0));

end fetchUnit;

architecture SYN_structural of fetchUnit is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component reg_12
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_0
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component IR
      port( clock, reset, load : in std_logic;  i : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux21_0
      port( a, b : in std_logic_vector (31 downto 0);  sel : in std_logic;  y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component Adder
      port( A, B : in std_logic_vector (31 downto 0);  reset, Cin : in 
            std_logic;  O : out std_logic_vector (31 downto 0);  Cout : out 
            std_logic);
   end component;
   
   signal X_Logic0_port, PCtoIM_31_port, PCtoIM_30_port, PCtoIM_29_port, 
      PCtoIM_28_port, PCtoIM_27_port, PCtoIM_26_port, PCtoIM_25_port, 
      PCtoIM_24_port, PCtoIM_23_port, PCtoIM_22_port, PCtoIM_21_port, 
      PCtoIM_20_port, PCtoIM_19_port, PCtoIM_18_port, PCtoIM_17_port, 
      PCtoIM_16_port, PCtoIM_15_port, PCtoIM_14_port, PCtoIM_13_port, 
      PCtoIM_12_port, PCtoIM_11_port, PCtoIM_10_port, PCtoIM_9_port, 
      PCtoIM_8_port, PCtoIM_7_port, PCtoIM_6_port, PCtoIM_5_port, PCtoIM_4_port
      , PCtoIM_3_port, PCtoIM_2_port, PCtoIM_1_port, PCtoIM_0_port, LOAD, 
      AddertoMux_31_port, AddertoMux_30_port, AddertoMux_29_port, 
      AddertoMux_28_port, AddertoMux_27_port, AddertoMux_26_port, 
      AddertoMux_25_port, AddertoMux_24_port, AddertoMux_23_port, 
      AddertoMux_22_port, AddertoMux_21_port, AddertoMux_20_port, 
      AddertoMux_19_port, AddertoMux_18_port, AddertoMux_17_port, 
      AddertoMux_16_port, AddertoMux_15_port, AddertoMux_14_port, 
      AddertoMux_13_port, AddertoMux_12_port, AddertoMux_11_port, 
      AddertoMux_10_port, AddertoMux_9_port, AddertoMux_8_port, 
      AddertoMux_7_port, AddertoMux_6_port, AddertoMux_5_port, 
      AddertoMux_4_port, AddertoMux_3_port, AddertoMux_2_port, 
      AddertoMux_1_port, AddertoMux_0_port, MuxtoPc_31_port, MuxtoPc_30_port, 
      MuxtoPc_29_port, MuxtoPc_28_port, MuxtoPc_27_port, MuxtoPc_26_port, 
      MuxtoPc_25_port, MuxtoPc_24_port, MuxtoPc_23_port, MuxtoPc_22_port, 
      MuxtoPc_21_port, MuxtoPc_20_port, MuxtoPc_19_port, MuxtoPc_18_port, 
      MuxtoPc_17_port, MuxtoPc_16_port, MuxtoPc_15_port, MuxtoPc_14_port, 
      MuxtoPc_13_port, MuxtoPc_12_port, MuxtoPc_11_port, MuxtoPc_10_port, 
      MuxtoPc_9_port, MuxtoPc_8_port, MuxtoPc_7_port, MuxtoPc_6_port, 
      MuxtoPc_5_port, MuxtoPc_4_port, MuxtoPc_3_port, MuxtoPc_2_port, 
      MuxtoPc_1_port, MuxtoPc_0_port, n_1353 : std_logic;

begin
   PCtoIM <= ( PCtoIM_31_port, PCtoIM_30_port, PCtoIM_29_port, PCtoIM_28_port, 
      PCtoIM_27_port, PCtoIM_26_port, PCtoIM_25_port, PCtoIM_24_port, 
      PCtoIM_23_port, PCtoIM_22_port, PCtoIM_21_port, PCtoIM_20_port, 
      PCtoIM_19_port, PCtoIM_18_port, PCtoIM_17_port, PCtoIM_16_port, 
      PCtoIM_15_port, PCtoIM_14_port, PCtoIM_13_port, PCtoIM_12_port, 
      PCtoIM_11_port, PCtoIM_10_port, PCtoIM_9_port, PCtoIM_8_port, 
      PCtoIM_7_port, PCtoIM_6_port, PCtoIM_5_port, PCtoIM_4_port, PCtoIM_3_port
      , PCtoIM_2_port, PCtoIM_1_port, PCtoIM_0_port );
   
   X_Logic0_port <= '0';
   nxpc : Adder port map( A(31) => PCtoIM_31_port, A(30) => PCtoIM_30_port, 
                           A(29) => PCtoIM_29_port, A(28) => PCtoIM_28_port, 
                           A(27) => PCtoIM_27_port, A(26) => PCtoIM_26_port, 
                           A(25) => PCtoIM_25_port, A(24) => PCtoIM_24_port, 
                           A(23) => PCtoIM_23_port, A(22) => PCtoIM_22_port, 
                           A(21) => PCtoIM_21_port, A(20) => PCtoIM_20_port, 
                           A(19) => PCtoIM_19_port, A(18) => PCtoIM_18_port, 
                           A(17) => PCtoIM_17_port, A(16) => PCtoIM_16_port, 
                           A(15) => PCtoIM_15_port, A(14) => PCtoIM_14_port, 
                           A(13) => PCtoIM_13_port, A(12) => PCtoIM_12_port, 
                           A(11) => PCtoIM_11_port, A(10) => PCtoIM_10_port, 
                           A(9) => PCtoIM_9_port, A(8) => PCtoIM_8_port, A(7) 
                           => PCtoIM_7_port, A(6) => PCtoIM_6_port, A(5) => 
                           PCtoIM_5_port, A(4) => PCtoIM_4_port, A(3) => 
                           PCtoIM_3_port, A(2) => PCtoIM_2_port, A(1) => 
                           PCtoIM_1_port, A(0) => PCtoIM_0_port, B(31) => 
                           X_Logic0_port, B(30) => X_Logic0_port, B(29) => 
                           X_Logic0_port, B(28) => X_Logic0_port, B(27) => 
                           X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
                           X_Logic0_port, B(24) => X_Logic0_port, B(23) => 
                           X_Logic0_port, B(22) => X_Logic0_port, B(21) => 
                           X_Logic0_port, B(20) => X_Logic0_port, B(19) => 
                           X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, reset => reset
                           , Cin => X_Logic0_port, O(31) => AddertoMux_31_port,
                           O(30) => AddertoMux_30_port, O(29) => 
                           AddertoMux_29_port, O(28) => AddertoMux_28_port, 
                           O(27) => AddertoMux_27_port, O(26) => 
                           AddertoMux_26_port, O(25) => AddertoMux_25_port, 
                           O(24) => AddertoMux_24_port, O(23) => 
                           AddertoMux_23_port, O(22) => AddertoMux_22_port, 
                           O(21) => AddertoMux_21_port, O(20) => 
                           AddertoMux_20_port, O(19) => AddertoMux_19_port, 
                           O(18) => AddertoMux_18_port, O(17) => 
                           AddertoMux_17_port, O(16) => AddertoMux_16_port, 
                           O(15) => AddertoMux_15_port, O(14) => 
                           AddertoMux_14_port, O(13) => AddertoMux_13_port, 
                           O(12) => AddertoMux_12_port, O(11) => 
                           AddertoMux_11_port, O(10) => AddertoMux_10_port, 
                           O(9) => AddertoMux_9_port, O(8) => AddertoMux_8_port
                           , O(7) => AddertoMux_7_port, O(6) => 
                           AddertoMux_6_port, O(5) => AddertoMux_5_port, O(4) 
                           => AddertoMux_4_port, O(3) => AddertoMux_3_port, 
                           O(2) => AddertoMux_2_port, O(1) => AddertoMux_1_port
                           , O(0) => AddertoMux_0_port, Cout => n_1353);
   pcmux : Mux21_0 port map( a(31) => BranchPC(31), a(30) => BranchPC(30), 
                           a(29) => BranchPC(29), a(28) => BranchPC(28), a(27) 
                           => BranchPC(27), a(26) => BranchPC(26), a(25) => 
                           BranchPC(25), a(24) => BranchPC(24), a(23) => 
                           BranchPC(23), a(22) => BranchPC(22), a(21) => 
                           BranchPC(21), a(20) => BranchPC(20), a(19) => 
                           BranchPC(19), a(18) => BranchPC(18), a(17) => 
                           BranchPC(17), a(16) => BranchPC(16), a(15) => 
                           BranchPC(15), a(14) => BranchPC(14), a(13) => 
                           BranchPC(13), a(12) => BranchPC(12), a(11) => 
                           BranchPC(11), a(10) => BranchPC(10), a(9) => 
                           BranchPC(9), a(8) => BranchPC(8), a(7) => 
                           BranchPC(7), a(6) => BranchPC(6), a(5) => 
                           BranchPC(5), a(4) => BranchPC(4), a(3) => 
                           BranchPC(3), a(2) => BranchPC(2), a(1) => 
                           BranchPC(1), a(0) => BranchPC(0), b(31) => 
                           AddertoMux_31_port, b(30) => AddertoMux_30_port, 
                           b(29) => AddertoMux_29_port, b(28) => 
                           AddertoMux_28_port, b(27) => AddertoMux_27_port, 
                           b(26) => AddertoMux_26_port, b(25) => 
                           AddertoMux_25_port, b(24) => AddertoMux_24_port, 
                           b(23) => AddertoMux_23_port, b(22) => 
                           AddertoMux_22_port, b(21) => AddertoMux_21_port, 
                           b(20) => AddertoMux_20_port, b(19) => 
                           AddertoMux_19_port, b(18) => AddertoMux_18_port, 
                           b(17) => AddertoMux_17_port, b(16) => 
                           AddertoMux_16_port, b(15) => AddertoMux_15_port, 
                           b(14) => AddertoMux_14_port, b(13) => 
                           AddertoMux_13_port, b(12) => AddertoMux_12_port, 
                           b(11) => AddertoMux_11_port, b(10) => 
                           AddertoMux_10_port, b(9) => AddertoMux_9_port, b(8) 
                           => AddertoMux_8_port, b(7) => AddertoMux_7_port, 
                           b(6) => AddertoMux_6_port, b(5) => AddertoMux_5_port
                           , b(4) => AddertoMux_4_port, b(3) => 
                           AddertoMux_3_port, b(2) => AddertoMux_2_port, b(1) 
                           => AddertoMux_1_port, b(0) => AddertoMux_0_port, sel
                           => BRANCHfromDECODE, y(31) => MuxtoPc_31_port, y(30)
                           => MuxtoPc_30_port, y(29) => MuxtoPc_29_port, y(28) 
                           => MuxtoPc_28_port, y(27) => MuxtoPc_27_port, y(26) 
                           => MuxtoPc_26_port, y(25) => MuxtoPc_25_port, y(24) 
                           => MuxtoPc_24_port, y(23) => MuxtoPc_23_port, y(22) 
                           => MuxtoPc_22_port, y(21) => MuxtoPc_21_port, y(20) 
                           => MuxtoPc_20_port, y(19) => MuxtoPc_19_port, y(18) 
                           => MuxtoPc_18_port, y(17) => MuxtoPc_17_port, y(16) 
                           => MuxtoPc_16_port, y(15) => MuxtoPc_15_port, y(14) 
                           => MuxtoPc_14_port, y(13) => MuxtoPc_13_port, y(12) 
                           => MuxtoPc_12_port, y(11) => MuxtoPc_11_port, y(10) 
                           => MuxtoPc_10_port, y(9) => MuxtoPc_9_port, y(8) => 
                           MuxtoPc_8_port, y(7) => MuxtoPc_7_port, y(6) => 
                           MuxtoPc_6_port, y(5) => MuxtoPc_5_port, y(4) => 
                           MuxtoPc_4_port, y(3) => MuxtoPc_3_port, y(2) => 
                           MuxtoPc_2_port, y(1) => MuxtoPc_1_port, y(0) => 
                           MuxtoPc_0_port);
   InstrReg : IR port map( clock => clock, reset => LOAD, load => en1, i(31) =>
                           Instruction(31), i(30) => Instruction(30), i(29) => 
                           Instruction(29), i(28) => Instruction(28), i(27) => 
                           Instruction(27), i(26) => Instruction(26), i(25) => 
                           Instruction(25), i(24) => Instruction(24), i(23) => 
                           Instruction(23), i(22) => Instruction(22), i(21) => 
                           Instruction(21), i(20) => Instruction(20), i(19) => 
                           Instruction(19), i(18) => Instruction(18), i(17) => 
                           Instruction(17), i(16) => Instruction(16), i(15) => 
                           Instruction(15), i(14) => Instruction(14), i(13) => 
                           Instruction(13), i(12) => Instruction(12), i(11) => 
                           Instruction(11), i(10) => Instruction(10), i(9) => 
                           Instruction(9), i(8) => Instruction(8), i(7) => 
                           Instruction(7), i(6) => Instruction(6), i(5) => 
                           Instruction(5), i(4) => Instruction(4), i(3) => 
                           Instruction(3), i(2) => Instruction(2), i(1) => 
                           Instruction(1), i(0) => Instruction(0), o(31) => 
                           IRtoDecode(31), o(30) => IRtoDecode(30), o(29) => 
                           IRtoDecode(29), o(28) => IRtoDecode(28), o(27) => 
                           IRtoDecode(27), o(26) => IRtoDecode(26), o(25) => 
                           IRtoDecode(25), o(24) => IRtoDecode(24), o(23) => 
                           IRtoDecode(23), o(22) => IRtoDecode(22), o(21) => 
                           IRtoDecode(21), o(20) => IRtoDecode(20), o(19) => 
                           IRtoDecode(19), o(18) => IRtoDecode(18), o(17) => 
                           IRtoDecode(17), o(16) => IRtoDecode(16), o(15) => 
                           IRtoDecode(15), o(14) => IRtoDecode(14), o(13) => 
                           IRtoDecode(13), o(12) => IRtoDecode(12), o(11) => 
                           IRtoDecode(11), o(10) => IRtoDecode(10), o(9) => 
                           IRtoDecode(9), o(8) => IRtoDecode(8), o(7) => 
                           IRtoDecode(7), o(6) => IRtoDecode(6), o(5) => 
                           IRtoDecode(5), o(4) => IRtoDecode(4), o(3) => 
                           IRtoDecode(3), o(2) => IRtoDecode(2), o(1) => 
                           IRtoDecode(1), o(0) => IRtoDecode(0));
   PC : reg_0 port map( clock => clock, reset => reset, load => en1, i(31) => 
                           MuxtoPc_31_port, i(30) => MuxtoPc_30_port, i(29) => 
                           MuxtoPc_29_port, i(28) => MuxtoPc_28_port, i(27) => 
                           MuxtoPc_27_port, i(26) => MuxtoPc_26_port, i(25) => 
                           MuxtoPc_25_port, i(24) => MuxtoPc_24_port, i(23) => 
                           MuxtoPc_23_port, i(22) => MuxtoPc_22_port, i(21) => 
                           MuxtoPc_21_port, i(20) => MuxtoPc_20_port, i(19) => 
                           MuxtoPc_19_port, i(18) => MuxtoPc_18_port, i(17) => 
                           MuxtoPc_17_port, i(16) => MuxtoPc_16_port, i(15) => 
                           MuxtoPc_15_port, i(14) => MuxtoPc_14_port, i(13) => 
                           MuxtoPc_13_port, i(12) => MuxtoPc_12_port, i(11) => 
                           MuxtoPc_11_port, i(10) => MuxtoPc_10_port, i(9) => 
                           MuxtoPc_9_port, i(8) => MuxtoPc_8_port, i(7) => 
                           MuxtoPc_7_port, i(6) => MuxtoPc_6_port, i(5) => 
                           MuxtoPc_5_port, i(4) => MuxtoPc_4_port, i(3) => 
                           MuxtoPc_3_port, i(2) => MuxtoPc_2_port, i(1) => 
                           MuxtoPc_1_port, i(0) => MuxtoPc_0_port, o(31) => 
                           PCtoIM_31_port, o(30) => PCtoIM_30_port, o(29) => 
                           PCtoIM_29_port, o(28) => PCtoIM_28_port, o(27) => 
                           PCtoIM_27_port, o(26) => PCtoIM_26_port, o(25) => 
                           PCtoIM_25_port, o(24) => PCtoIM_24_port, o(23) => 
                           PCtoIM_23_port, o(22) => PCtoIM_22_port, o(21) => 
                           PCtoIM_21_port, o(20) => PCtoIM_20_port, o(19) => 
                           PCtoIM_19_port, o(18) => PCtoIM_18_port, o(17) => 
                           PCtoIM_17_port, o(16) => PCtoIM_16_port, o(15) => 
                           PCtoIM_15_port, o(14) => PCtoIM_14_port, o(13) => 
                           PCtoIM_13_port, o(12) => PCtoIM_12_port, o(11) => 
                           PCtoIM_11_port, o(10) => PCtoIM_10_port, o(9) => 
                           PCtoIM_9_port, o(8) => PCtoIM_8_port, o(7) => 
                           PCtoIM_7_port, o(6) => PCtoIM_6_port, o(5) => 
                           PCtoIM_5_port, o(4) => PCtoIM_4_port, o(3) => 
                           PCtoIM_3_port, o(2) => PCtoIM_2_port, o(1) => 
                           PCtoIM_1_port, o(0) => PCtoIM_0_port);
   NPC : reg_12 port map( clock => clock, reset => reset, load => en1, i(31) =>
                           AddertoMux_31_port, i(30) => AddertoMux_30_port, 
                           i(29) => AddertoMux_29_port, i(28) => 
                           AddertoMux_28_port, i(27) => AddertoMux_27_port, 
                           i(26) => AddertoMux_26_port, i(25) => 
                           AddertoMux_25_port, i(24) => AddertoMux_24_port, 
                           i(23) => AddertoMux_23_port, i(22) => 
                           AddertoMux_22_port, i(21) => AddertoMux_21_port, 
                           i(20) => AddertoMux_20_port, i(19) => 
                           AddertoMux_19_port, i(18) => AddertoMux_18_port, 
                           i(17) => AddertoMux_17_port, i(16) => 
                           AddertoMux_16_port, i(15) => AddertoMux_15_port, 
                           i(14) => AddertoMux_14_port, i(13) => 
                           AddertoMux_13_port, i(12) => AddertoMux_12_port, 
                           i(11) => AddertoMux_11_port, i(10) => 
                           AddertoMux_10_port, i(9) => AddertoMux_9_port, i(8) 
                           => AddertoMux_8_port, i(7) => AddertoMux_7_port, 
                           i(6) => AddertoMux_6_port, i(5) => AddertoMux_5_port
                           , i(4) => AddertoMux_4_port, i(3) => 
                           AddertoMux_3_port, i(2) => AddertoMux_2_port, i(1) 
                           => AddertoMux_1_port, i(0) => AddertoMux_0_port, 
                           o(31) => NPCtoDecode(31), o(30) => NPCtoDecode(30), 
                           o(29) => NPCtoDecode(29), o(28) => NPCtoDecode(28), 
                           o(27) => NPCtoDecode(27), o(26) => NPCtoDecode(26), 
                           o(25) => NPCtoDecode(25), o(24) => NPCtoDecode(24), 
                           o(23) => NPCtoDecode(23), o(22) => NPCtoDecode(22), 
                           o(21) => NPCtoDecode(21), o(20) => NPCtoDecode(20), 
                           o(19) => NPCtoDecode(19), o(18) => NPCtoDecode(18), 
                           o(17) => NPCtoDecode(17), o(16) => NPCtoDecode(16), 
                           o(15) => NPCtoDecode(15), o(14) => NPCtoDecode(14), 
                           o(13) => NPCtoDecode(13), o(12) => NPCtoDecode(12), 
                           o(11) => NPCtoDecode(11), o(10) => NPCtoDecode(10), 
                           o(9) => NPCtoDecode(9), o(8) => NPCtoDecode(8), o(7)
                           => NPCtoDecode(7), o(6) => NPCtoDecode(6), o(5) => 
                           NPCtoDecode(5), o(4) => NPCtoDecode(4), o(3) => 
                           NPCtoDecode(3), o(2) => NPCtoDecode(2), o(1) => 
                           NPCtoDecode(1), o(0) => NPCtoDecode(0));
   U2 : OR2_X1 port map( A1 => BRANCHfromDECODE, A2 => reset, ZN => LOAD);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity dataPath_M32_C4_N5 is

   port( clock, reset : in std_logic;  Instruction : in std_logic_vector (31 
         downto 0);  en1, en2, SignSelect, RD1, RD2, WR, JMP, BRANCHenable, en3
         , BranchCondSel, Mux1Sel, Mux2Sel : in std_logic;  ALUCODE : in 
         std_logic_vector (3 downto 0);  RegDestination, en4 : in std_logic;  
         DRAMout : in std_logic_vector (31 downto 0);  selwb : in std_logic;  
         PCtoIM, ALUtoMEMORY, OUT2RFtoMEMORY, InstructionToCU : out 
         std_logic_vector (31 downto 0));

end dataPath_M32_C4_N5;

architecture SYN_structural of dataPath_M32_C4_N5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component WBUnit
      port( selwb : in std_logic;  ALUin, LOADDATA, AddressWfromMemory : in 
            std_logic_vector (31 downto 0);  MUXtoRF, AddressWtoDECODE : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component memoryUnit
      port( clock, reset, en4 : in std_logic;  ALUout, DRAMout, 
            AddressWfromEXECUTE : in std_logic_vector (31 downto 0);  LOADDATA,
            ALUtoWBMUX, AddressWtoWB : out std_logic_vector (31 downto 0));
   end component;
   
   component executeUnit_M32_C4
      port( clock, reset, en3, Mux1Sel, Mux2Sel : in std_logic;  ALUCODE : in 
            std_logic_vector (3 downto 0);  OUT1RF, OUT2RF, IMMEDIATE, 
            NPCFromDecode, AddressWfromDecode : in std_logic_vector (31 downto 
            0);  ALUtoMEMORY, OUT2RFtoMEMORY, AddressWtoMEMORY : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component DecodeUnit
      port( clock, reset, JMP, RegDestination, en2, SignSelect, BranchCondSel, 
            BRANCHenable, RD1, RD2, WR : in std_logic;  Instruction : in 
            std_logic_vector (31 downto 0);  ADD_WR : in std_logic_vector (4 
            downto 0);  DATAIN, NPCfromIF : in std_logic_vector (31 downto 0); 
            OUT1, OUT2, OUTNPC, OUTIMM, NPCtoEX, AddressWtoEX : out 
            std_logic_vector (31 downto 0);  BRANCHtoFetch : out std_logic);
   end component;
   
   component fetchUnit
      port( clock, reset, en1 : in std_logic;  BranchPC : in std_logic_vector 
            (31 downto 0);  BRANCHfromDECODE : in std_logic;  Instruction : in 
            std_logic_vector (31 downto 0);  PCtoIM, IRtoDecode, NPCtoDecode : 
            out std_logic_vector (31 downto 0));
   end component;
   
   signal ALUtoMEMORY_31_port, ALUtoMEMORY_30_port, ALUtoMEMORY_29_port, 
      ALUtoMEMORY_28_port, ALUtoMEMORY_27_port, ALUtoMEMORY_26_port, 
      ALUtoMEMORY_25_port, ALUtoMEMORY_24_port, ALUtoMEMORY_23_port, 
      ALUtoMEMORY_22_port, ALUtoMEMORY_21_port, ALUtoMEMORY_20_port, 
      ALUtoMEMORY_19_port, ALUtoMEMORY_18_port, ALUtoMEMORY_17_port, 
      ALUtoMEMORY_16_port, ALUtoMEMORY_15_port, ALUtoMEMORY_14_port, 
      ALUtoMEMORY_13_port, ALUtoMEMORY_12_port, ALUtoMEMORY_11_port, 
      ALUtoMEMORY_10_port, ALUtoMEMORY_9_port, ALUtoMEMORY_8_port, 
      ALUtoMEMORY_7_port, ALUtoMEMORY_6_port, ALUtoMEMORY_5_port, 
      ALUtoMEMORY_4_port, ALUtoMEMORY_3_port, ALUtoMEMORY_2_port, 
      ALUtoMEMORY_1_port, ALUtoMEMORY_0_port, InstructionToCU_31_port, 
      InstructionToCU_30_port, InstructionToCU_29_port, InstructionToCU_28_port
      , InstructionToCU_27_port, InstructionToCU_26_port, 
      InstructionToCU_25_port, InstructionToCU_24_port, InstructionToCU_23_port
      , InstructionToCU_22_port, InstructionToCU_21_port, 
      InstructionToCU_20_port, InstructionToCU_19_port, InstructionToCU_18_port
      , InstructionToCU_17_port, InstructionToCU_16_port, 
      InstructionToCU_15_port, InstructionToCU_14_port, InstructionToCU_13_port
      , InstructionToCU_12_port, InstructionToCU_11_port, 
      InstructionToCU_10_port, InstructionToCU_9_port, InstructionToCU_8_port, 
      InstructionToCU_7_port, InstructionToCU_6_port, InstructionToCU_5_port, 
      InstructionToCU_4_port, InstructionToCU_3_port, InstructionToCU_2_port, 
      InstructionToCU_1_port, InstructionToCU_0_port, NewPC_31_port, 
      NewPC_30_port, NewPC_29_port, NewPC_28_port, NewPC_27_port, NewPC_26_port
      , NewPC_25_port, NewPC_24_port, NewPC_23_port, NewPC_22_port, 
      NewPC_21_port, NewPC_20_port, NewPC_19_port, NewPC_18_port, NewPC_17_port
      , NewPC_16_port, NewPC_15_port, NewPC_14_port, NewPC_13_port, 
      NewPC_12_port, NewPC_11_port, NewPC_10_port, NewPC_9_port, NewPC_8_port, 
      NewPC_7_port, NewPC_6_port, NewPC_5_port, NewPC_4_port, NewPC_3_port, 
      NewPC_2_port, NewPC_1_port, NewPC_0_port, BRANCHtoFetch, NXPC_31_port, 
      NXPC_30_port, NXPC_29_port, NXPC_28_port, NXPC_27_port, NXPC_26_port, 
      NXPC_25_port, NXPC_24_port, NXPC_23_port, NXPC_22_port, NXPC_21_port, 
      NXPC_20_port, NXPC_19_port, NXPC_18_port, NXPC_17_port, NXPC_16_port, 
      NXPC_15_port, NXPC_14_port, NXPC_13_port, NXPC_12_port, NXPC_11_port, 
      NXPC_10_port, NXPC_9_port, NXPC_8_port, NXPC_7_port, NXPC_6_port, 
      NXPC_5_port, NXPC_4_port, NXPC_3_port, NXPC_2_port, NXPC_1_port, 
      NXPC_0_port, AddressfromWB_4_port, AddressfromWB_3_port, 
      AddressfromWB_2_port, AddressfromWB_1_port, AddressfromWB_0_port, 
      MUXtoRF_31_port, MUXtoRF_30_port, MUXtoRF_29_port, MUXtoRF_28_port, 
      MUXtoRF_27_port, MUXtoRF_26_port, MUXtoRF_25_port, MUXtoRF_24_port, 
      MUXtoRF_23_port, MUXtoRF_22_port, MUXtoRF_21_port, MUXtoRF_20_port, 
      MUXtoRF_19_port, MUXtoRF_18_port, MUXtoRF_17_port, MUXtoRF_16_port, 
      MUXtoRF_15_port, MUXtoRF_14_port, MUXtoRF_13_port, MUXtoRF_12_port, 
      MUXtoRF_11_port, MUXtoRF_10_port, MUXtoRF_9_port, MUXtoRF_8_port, 
      MUXtoRF_7_port, MUXtoRF_6_port, MUXtoRF_5_port, MUXtoRF_4_port, 
      MUXtoRF_3_port, MUXtoRF_2_port, MUXtoRF_1_port, MUXtoRF_0_port, 
      OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port, 
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, 
      OUT1_1_port, OUT1_0_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, 
      OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, 
      OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, 
      OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, 
      OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, 
      OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, 
      OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port, OUTIMM_31_port, 
      OUTIMM_30_port, OUTIMM_29_port, OUTIMM_28_port, OUTIMM_27_port, 
      OUTIMM_26_port, OUTIMM_25_port, OUTIMM_24_port, OUTIMM_23_port, 
      OUTIMM_22_port, OUTIMM_21_port, OUTIMM_20_port, OUTIMM_19_port, 
      OUTIMM_18_port, OUTIMM_17_port, OUTIMM_16_port, OUTIMM_15_port, 
      OUTIMM_14_port, OUTIMM_13_port, OUTIMM_12_port, OUTIMM_11_port, 
      OUTIMM_10_port, OUTIMM_9_port, OUTIMM_8_port, OUTIMM_7_port, 
      OUTIMM_6_port, OUTIMM_5_port, OUTIMM_4_port, OUTIMM_3_port, OUTIMM_2_port
      , OUTIMM_1_port, OUTIMM_0_port, NPCfromDECODE_31_port, 
      NPCfromDECODE_30_port, NPCfromDECODE_29_port, NPCfromDECODE_28_port, 
      NPCfromDECODE_27_port, NPCfromDECODE_26_port, NPCfromDECODE_25_port, 
      NPCfromDECODE_24_port, NPCfromDECODE_23_port, NPCfromDECODE_22_port, 
      NPCfromDECODE_21_port, NPCfromDECODE_20_port, NPCfromDECODE_19_port, 
      NPCfromDECODE_18_port, NPCfromDECODE_17_port, NPCfromDECODE_16_port, 
      NPCfromDECODE_15_port, NPCfromDECODE_14_port, NPCfromDECODE_13_port, 
      NPCfromDECODE_12_port, NPCfromDECODE_11_port, NPCfromDECODE_10_port, 
      NPCfromDECODE_9_port, NPCfromDECODE_8_port, NPCfromDECODE_7_port, 
      NPCfromDECODE_6_port, NPCfromDECODE_5_port, NPCfromDECODE_4_port, 
      NPCfromDECODE_3_port, NPCfromDECODE_2_port, NPCfromDECODE_1_port, 
      NPCfromDECODE_0_port, ADDWfromDECODE_31_port, ADDWfromDECODE_30_port, 
      ADDWfromDECODE_29_port, ADDWfromDECODE_28_port, ADDWfromDECODE_27_port, 
      ADDWfromDECODE_26_port, ADDWfromDECODE_25_port, ADDWfromDECODE_24_port, 
      ADDWfromDECODE_23_port, ADDWfromDECODE_22_port, ADDWfromDECODE_21_port, 
      ADDWfromDECODE_20_port, ADDWfromDECODE_19_port, ADDWfromDECODE_18_port, 
      ADDWfromDECODE_17_port, ADDWfromDECODE_16_port, ADDWfromDECODE_15_port, 
      ADDWfromDECODE_14_port, ADDWfromDECODE_13_port, ADDWfromDECODE_12_port, 
      ADDWfromDECODE_11_port, ADDWfromDECODE_10_port, ADDWfromDECODE_9_port, 
      ADDWfromDECODE_8_port, ADDWfromDECODE_7_port, ADDWfromDECODE_6_port, 
      ADDWfromDECODE_5_port, ADDWfromDECODE_4_port, ADDWfromDECODE_3_port, 
      ADDWfromDECODE_2_port, ADDWfromDECODE_1_port, ADDWfromDECODE_0_port, 
      ADDWtoMEMORY_31_port, ADDWtoMEMORY_30_port, ADDWtoMEMORY_29_port, 
      ADDWtoMEMORY_28_port, ADDWtoMEMORY_27_port, ADDWtoMEMORY_26_port, 
      ADDWtoMEMORY_25_port, ADDWtoMEMORY_24_port, ADDWtoMEMORY_23_port, 
      ADDWtoMEMORY_22_port, ADDWtoMEMORY_21_port, ADDWtoMEMORY_20_port, 
      ADDWtoMEMORY_19_port, ADDWtoMEMORY_18_port, ADDWtoMEMORY_17_port, 
      ADDWtoMEMORY_16_port, ADDWtoMEMORY_15_port, ADDWtoMEMORY_14_port, 
      ADDWtoMEMORY_13_port, ADDWtoMEMORY_12_port, ADDWtoMEMORY_11_port, 
      ADDWtoMEMORY_10_port, ADDWtoMEMORY_9_port, ADDWtoMEMORY_8_port, 
      ADDWtoMEMORY_7_port, ADDWtoMEMORY_6_port, ADDWtoMEMORY_5_port, 
      ADDWtoMEMORY_4_port, ADDWtoMEMORY_3_port, ADDWtoMEMORY_2_port, 
      ADDWtoMEMORY_1_port, ADDWtoMEMORY_0_port, LOADDATA_31_port, 
      LOADDATA_30_port, LOADDATA_29_port, LOADDATA_28_port, LOADDATA_27_port, 
      LOADDATA_26_port, LOADDATA_25_port, LOADDATA_24_port, LOADDATA_23_port, 
      LOADDATA_22_port, LOADDATA_21_port, LOADDATA_20_port, LOADDATA_19_port, 
      LOADDATA_18_port, LOADDATA_17_port, LOADDATA_16_port, LOADDATA_15_port, 
      LOADDATA_14_port, LOADDATA_13_port, LOADDATA_12_port, LOADDATA_11_port, 
      LOADDATA_10_port, LOADDATA_9_port, LOADDATA_8_port, LOADDATA_7_port, 
      LOADDATA_6_port, LOADDATA_5_port, LOADDATA_4_port, LOADDATA_3_port, 
      LOADDATA_2_port, LOADDATA_1_port, LOADDATA_0_port, ALUtoWBMUX_31_port, 
      ALUtoWBMUX_30_port, ALUtoWBMUX_29_port, ALUtoWBMUX_28_port, 
      ALUtoWBMUX_27_port, ALUtoWBMUX_26_port, ALUtoWBMUX_25_port, 
      ALUtoWBMUX_24_port, ALUtoWBMUX_23_port, ALUtoWBMUX_22_port, 
      ALUtoWBMUX_21_port, ALUtoWBMUX_20_port, ALUtoWBMUX_19_port, 
      ALUtoWBMUX_18_port, ALUtoWBMUX_17_port, ALUtoWBMUX_16_port, 
      ALUtoWBMUX_15_port, ALUtoWBMUX_14_port, ALUtoWBMUX_13_port, 
      ALUtoWBMUX_12_port, ALUtoWBMUX_11_port, ALUtoWBMUX_10_port, 
      ALUtoWBMUX_9_port, ALUtoWBMUX_8_port, ALUtoWBMUX_7_port, 
      ALUtoWBMUX_6_port, ALUtoWBMUX_5_port, ALUtoWBMUX_4_port, 
      ALUtoWBMUX_3_port, ALUtoWBMUX_2_port, ALUtoWBMUX_1_port, 
      ALUtoWBMUX_0_port, ADDWtoWB_31_port, ADDWtoWB_30_port, ADDWtoWB_29_port, 
      ADDWtoWB_28_port, ADDWtoWB_27_port, ADDWtoWB_26_port, ADDWtoWB_25_port, 
      ADDWtoWB_24_port, ADDWtoWB_23_port, ADDWtoWB_22_port, ADDWtoWB_21_port, 
      ADDWtoWB_20_port, ADDWtoWB_19_port, ADDWtoWB_18_port, ADDWtoWB_17_port, 
      ADDWtoWB_16_port, ADDWtoWB_15_port, ADDWtoWB_14_port, ADDWtoWB_13_port, 
      ADDWtoWB_12_port, ADDWtoWB_11_port, ADDWtoWB_10_port, ADDWtoWB_9_port, 
      ADDWtoWB_8_port, ADDWtoWB_7_port, ADDWtoWB_6_port, ADDWtoWB_5_port, 
      ADDWtoWB_4_port, ADDWtoWB_3_port, ADDWtoWB_2_port, ADDWtoWB_1_port, 
      ADDWtoWB_0_port, n1, n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, 
      n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, 
      n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, 
      n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, 
      n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, 
      n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402 : std_logic;

begin
   ALUtoMEMORY <= ( ALUtoMEMORY_31_port, ALUtoMEMORY_30_port, 
      ALUtoMEMORY_29_port, ALUtoMEMORY_28_port, ALUtoMEMORY_27_port, 
      ALUtoMEMORY_26_port, ALUtoMEMORY_25_port, ALUtoMEMORY_24_port, 
      ALUtoMEMORY_23_port, ALUtoMEMORY_22_port, ALUtoMEMORY_21_port, 
      ALUtoMEMORY_20_port, ALUtoMEMORY_19_port, ALUtoMEMORY_18_port, 
      ALUtoMEMORY_17_port, ALUtoMEMORY_16_port, ALUtoMEMORY_15_port, 
      ALUtoMEMORY_14_port, ALUtoMEMORY_13_port, ALUtoMEMORY_12_port, 
      ALUtoMEMORY_11_port, ALUtoMEMORY_10_port, ALUtoMEMORY_9_port, 
      ALUtoMEMORY_8_port, ALUtoMEMORY_7_port, ALUtoMEMORY_6_port, 
      ALUtoMEMORY_5_port, ALUtoMEMORY_4_port, ALUtoMEMORY_3_port, 
      ALUtoMEMORY_2_port, ALUtoMEMORY_1_port, ALUtoMEMORY_0_port );
   InstructionToCU <= ( InstructionToCU_31_port, InstructionToCU_30_port, 
      InstructionToCU_29_port, InstructionToCU_28_port, InstructionToCU_27_port
      , InstructionToCU_26_port, InstructionToCU_25_port, 
      InstructionToCU_24_port, InstructionToCU_23_port, InstructionToCU_22_port
      , InstructionToCU_21_port, InstructionToCU_20_port, 
      InstructionToCU_19_port, InstructionToCU_18_port, InstructionToCU_17_port
      , InstructionToCU_16_port, InstructionToCU_15_port, 
      InstructionToCU_14_port, InstructionToCU_13_port, InstructionToCU_12_port
      , InstructionToCU_11_port, InstructionToCU_10_port, 
      InstructionToCU_9_port, InstructionToCU_8_port, InstructionToCU_7_port, 
      InstructionToCU_6_port, InstructionToCU_5_port, InstructionToCU_4_port, 
      InstructionToCU_3_port, InstructionToCU_2_port, InstructionToCU_1_port, 
      InstructionToCU_0_port );
   
   NewPC_10_port <= '0';
   NewPC_11_port <= '0';
   NewPC_12_port <= '0';
   NewPC_13_port <= '0';
   NewPC_14_port <= '0';
   NewPC_15_port <= '0';
   NewPC_16_port <= '0';
   NewPC_17_port <= '0';
   NewPC_18_port <= '0';
   NewPC_19_port <= '0';
   NewPC_20_port <= '0';
   NewPC_21_port <= '0';
   NewPC_22_port <= '0';
   NewPC_23_port <= '0';
   NewPC_24_port <= '0';
   NewPC_25_port <= '0';
   NewPC_26_port <= '0';
   NewPC_27_port <= '0';
   NewPC_28_port <= '0';
   NewPC_29_port <= '0';
   NewPC_30_port <= '0';
   NewPC_31_port <= '0';
   FU : fetchUnit port map( clock => clock, reset => n1, en1 => en1, 
                           BranchPC(31) => NewPC_31_port, BranchPC(30) => 
                           NewPC_30_port, BranchPC(29) => NewPC_29_port, 
                           BranchPC(28) => NewPC_28_port, BranchPC(27) => 
                           NewPC_27_port, BranchPC(26) => NewPC_26_port, 
                           BranchPC(25) => NewPC_25_port, BranchPC(24) => 
                           NewPC_24_port, BranchPC(23) => NewPC_23_port, 
                           BranchPC(22) => NewPC_22_port, BranchPC(21) => 
                           NewPC_21_port, BranchPC(20) => NewPC_20_port, 
                           BranchPC(19) => NewPC_19_port, BranchPC(18) => 
                           NewPC_18_port, BranchPC(17) => NewPC_17_port, 
                           BranchPC(16) => NewPC_16_port, BranchPC(15) => 
                           NewPC_15_port, BranchPC(14) => NewPC_14_port, 
                           BranchPC(13) => NewPC_13_port, BranchPC(12) => 
                           NewPC_12_port, BranchPC(11) => NewPC_11_port, 
                           BranchPC(10) => NewPC_10_port, BranchPC(9) => 
                           NewPC_9_port, BranchPC(8) => NewPC_8_port, 
                           BranchPC(7) => NewPC_7_port, BranchPC(6) => 
                           NewPC_6_port, BranchPC(5) => NewPC_5_port, 
                           BranchPC(4) => NewPC_4_port, BranchPC(3) => 
                           NewPC_3_port, BranchPC(2) => NewPC_2_port, 
                           BranchPC(1) => NewPC_1_port, BranchPC(0) => 
                           NewPC_0_port, BRANCHfromDECODE => BRANCHtoFetch, 
                           Instruction(31) => Instruction(31), Instruction(30) 
                           => Instruction(30), Instruction(29) => 
                           Instruction(29), Instruction(28) => Instruction(28),
                           Instruction(27) => Instruction(27), Instruction(26) 
                           => Instruction(26), Instruction(25) => 
                           Instruction(25), Instruction(24) => Instruction(24),
                           Instruction(23) => Instruction(23), Instruction(22) 
                           => Instruction(22), Instruction(21) => 
                           Instruction(21), Instruction(20) => Instruction(20),
                           Instruction(19) => Instruction(19), Instruction(18) 
                           => Instruction(18), Instruction(17) => 
                           Instruction(17), Instruction(16) => Instruction(16),
                           Instruction(15) => Instruction(15), Instruction(14) 
                           => Instruction(14), Instruction(13) => 
                           Instruction(13), Instruction(12) => Instruction(12),
                           Instruction(11) => Instruction(11), Instruction(10) 
                           => Instruction(10), Instruction(9) => Instruction(9)
                           , Instruction(8) => Instruction(8), Instruction(7) 
                           => Instruction(7), Instruction(6) => Instruction(6),
                           Instruction(5) => Instruction(5), Instruction(4) => 
                           Instruction(4), Instruction(3) => Instruction(3), 
                           Instruction(2) => Instruction(2), Instruction(1) => 
                           Instruction(1), Instruction(0) => Instruction(0), 
                           PCtoIM(31) => PCtoIM(31), PCtoIM(30) => PCtoIM(30), 
                           PCtoIM(29) => PCtoIM(29), PCtoIM(28) => PCtoIM(28), 
                           PCtoIM(27) => PCtoIM(27), PCtoIM(26) => PCtoIM(26), 
                           PCtoIM(25) => PCtoIM(25), PCtoIM(24) => PCtoIM(24), 
                           PCtoIM(23) => PCtoIM(23), PCtoIM(22) => PCtoIM(22), 
                           PCtoIM(21) => PCtoIM(21), PCtoIM(20) => PCtoIM(20), 
                           PCtoIM(19) => PCtoIM(19), PCtoIM(18) => PCtoIM(18), 
                           PCtoIM(17) => PCtoIM(17), PCtoIM(16) => PCtoIM(16), 
                           PCtoIM(15) => PCtoIM(15), PCtoIM(14) => PCtoIM(14), 
                           PCtoIM(13) => PCtoIM(13), PCtoIM(12) => PCtoIM(12), 
                           PCtoIM(11) => PCtoIM(11), PCtoIM(10) => PCtoIM(10), 
                           PCtoIM(9) => PCtoIM(9), PCtoIM(8) => PCtoIM(8), 
                           PCtoIM(7) => PCtoIM(7), PCtoIM(6) => PCtoIM(6), 
                           PCtoIM(5) => PCtoIM(5), PCtoIM(4) => PCtoIM(4), 
                           PCtoIM(3) => PCtoIM(3), PCtoIM(2) => PCtoIM(2), 
                           PCtoIM(1) => PCtoIM(1), PCtoIM(0) => PCtoIM(0), 
                           IRtoDecode(31) => InstructionToCU_31_port, 
                           IRtoDecode(30) => InstructionToCU_30_port, 
                           IRtoDecode(29) => InstructionToCU_29_port, 
                           IRtoDecode(28) => InstructionToCU_28_port, 
                           IRtoDecode(27) => InstructionToCU_27_port, 
                           IRtoDecode(26) => InstructionToCU_26_port, 
                           IRtoDecode(25) => InstructionToCU_25_port, 
                           IRtoDecode(24) => InstructionToCU_24_port, 
                           IRtoDecode(23) => InstructionToCU_23_port, 
                           IRtoDecode(22) => InstructionToCU_22_port, 
                           IRtoDecode(21) => InstructionToCU_21_port, 
                           IRtoDecode(20) => InstructionToCU_20_port, 
                           IRtoDecode(19) => InstructionToCU_19_port, 
                           IRtoDecode(18) => InstructionToCU_18_port, 
                           IRtoDecode(17) => InstructionToCU_17_port, 
                           IRtoDecode(16) => InstructionToCU_16_port, 
                           IRtoDecode(15) => InstructionToCU_15_port, 
                           IRtoDecode(14) => InstructionToCU_14_port, 
                           IRtoDecode(13) => InstructionToCU_13_port, 
                           IRtoDecode(12) => InstructionToCU_12_port, 
                           IRtoDecode(11) => InstructionToCU_11_port, 
                           IRtoDecode(10) => InstructionToCU_10_port, 
                           IRtoDecode(9) => InstructionToCU_9_port, 
                           IRtoDecode(8) => InstructionToCU_8_port, 
                           IRtoDecode(7) => InstructionToCU_7_port, 
                           IRtoDecode(6) => InstructionToCU_6_port, 
                           IRtoDecode(5) => InstructionToCU_5_port, 
                           IRtoDecode(4) => InstructionToCU_4_port, 
                           IRtoDecode(3) => InstructionToCU_3_port, 
                           IRtoDecode(2) => InstructionToCU_2_port, 
                           IRtoDecode(1) => InstructionToCU_1_port, 
                           IRtoDecode(0) => InstructionToCU_0_port, 
                           NPCtoDecode(31) => NXPC_31_port, NPCtoDecode(30) => 
                           NXPC_30_port, NPCtoDecode(29) => NXPC_29_port, 
                           NPCtoDecode(28) => NXPC_28_port, NPCtoDecode(27) => 
                           NXPC_27_port, NPCtoDecode(26) => NXPC_26_port, 
                           NPCtoDecode(25) => NXPC_25_port, NPCtoDecode(24) => 
                           NXPC_24_port, NPCtoDecode(23) => NXPC_23_port, 
                           NPCtoDecode(22) => NXPC_22_port, NPCtoDecode(21) => 
                           NXPC_21_port, NPCtoDecode(20) => NXPC_20_port, 
                           NPCtoDecode(19) => NXPC_19_port, NPCtoDecode(18) => 
                           NXPC_18_port, NPCtoDecode(17) => NXPC_17_port, 
                           NPCtoDecode(16) => NXPC_16_port, NPCtoDecode(15) => 
                           NXPC_15_port, NPCtoDecode(14) => NXPC_14_port, 
                           NPCtoDecode(13) => NXPC_13_port, NPCtoDecode(12) => 
                           NXPC_12_port, NPCtoDecode(11) => NXPC_11_port, 
                           NPCtoDecode(10) => NXPC_10_port, NPCtoDecode(9) => 
                           NXPC_9_port, NPCtoDecode(8) => NXPC_8_port, 
                           NPCtoDecode(7) => NXPC_7_port, NPCtoDecode(6) => 
                           NXPC_6_port, NPCtoDecode(5) => NXPC_5_port, 
                           NPCtoDecode(4) => NXPC_4_port, NPCtoDecode(3) => 
                           NXPC_3_port, NPCtoDecode(2) => NXPC_2_port, 
                           NPCtoDecode(1) => NXPC_1_port, NPCtoDecode(0) => 
                           NXPC_0_port);
   DU : DecodeUnit port map( clock => clock, reset => n1, JMP => JMP, 
                           RegDestination => RegDestination, en2 => en2, 
                           SignSelect => SignSelect, BranchCondSel => 
                           BranchCondSel, BRANCHenable => BRANCHenable, RD1 => 
                           RD1, RD2 => RD2, WR => WR, Instruction(31) => 
                           InstructionToCU_31_port, Instruction(30) => 
                           InstructionToCU_30_port, Instruction(29) => 
                           InstructionToCU_29_port, Instruction(28) => 
                           InstructionToCU_28_port, Instruction(27) => 
                           InstructionToCU_27_port, Instruction(26) => 
                           InstructionToCU_26_port, Instruction(25) => 
                           InstructionToCU_25_port, Instruction(24) => 
                           InstructionToCU_24_port, Instruction(23) => 
                           InstructionToCU_23_port, Instruction(22) => 
                           InstructionToCU_22_port, Instruction(21) => 
                           InstructionToCU_21_port, Instruction(20) => 
                           InstructionToCU_20_port, Instruction(19) => 
                           InstructionToCU_19_port, Instruction(18) => 
                           InstructionToCU_18_port, Instruction(17) => 
                           InstructionToCU_17_port, Instruction(16) => 
                           InstructionToCU_16_port, Instruction(15) => 
                           InstructionToCU_15_port, Instruction(14) => 
                           InstructionToCU_14_port, Instruction(13) => 
                           InstructionToCU_13_port, Instruction(12) => 
                           InstructionToCU_12_port, Instruction(11) => 
                           InstructionToCU_11_port, Instruction(10) => 
                           InstructionToCU_10_port, Instruction(9) => 
                           InstructionToCU_9_port, Instruction(8) => 
                           InstructionToCU_8_port, Instruction(7) => 
                           InstructionToCU_7_port, Instruction(6) => 
                           InstructionToCU_6_port, Instruction(5) => 
                           InstructionToCU_5_port, Instruction(4) => 
                           InstructionToCU_4_port, Instruction(3) => 
                           InstructionToCU_3_port, Instruction(2) => 
                           InstructionToCU_2_port, Instruction(1) => 
                           InstructionToCU_1_port, Instruction(0) => 
                           InstructionToCU_0_port, ADD_WR(4) => 
                           AddressfromWB_4_port, ADD_WR(3) => 
                           AddressfromWB_3_port, ADD_WR(2) => 
                           AddressfromWB_2_port, ADD_WR(1) => 
                           AddressfromWB_1_port, ADD_WR(0) => 
                           AddressfromWB_0_port, DATAIN(31) => MUXtoRF_31_port,
                           DATAIN(30) => MUXtoRF_30_port, DATAIN(29) => 
                           MUXtoRF_29_port, DATAIN(28) => MUXtoRF_28_port, 
                           DATAIN(27) => MUXtoRF_27_port, DATAIN(26) => 
                           MUXtoRF_26_port, DATAIN(25) => MUXtoRF_25_port, 
                           DATAIN(24) => MUXtoRF_24_port, DATAIN(23) => 
                           MUXtoRF_23_port, DATAIN(22) => MUXtoRF_22_port, 
                           DATAIN(21) => MUXtoRF_21_port, DATAIN(20) => 
                           MUXtoRF_20_port, DATAIN(19) => MUXtoRF_19_port, 
                           DATAIN(18) => MUXtoRF_18_port, DATAIN(17) => 
                           MUXtoRF_17_port, DATAIN(16) => MUXtoRF_16_port, 
                           DATAIN(15) => MUXtoRF_15_port, DATAIN(14) => 
                           MUXtoRF_14_port, DATAIN(13) => MUXtoRF_13_port, 
                           DATAIN(12) => MUXtoRF_12_port, DATAIN(11) => 
                           MUXtoRF_11_port, DATAIN(10) => MUXtoRF_10_port, 
                           DATAIN(9) => MUXtoRF_9_port, DATAIN(8) => 
                           MUXtoRF_8_port, DATAIN(7) => MUXtoRF_7_port, 
                           DATAIN(6) => MUXtoRF_6_port, DATAIN(5) => 
                           MUXtoRF_5_port, DATAIN(4) => MUXtoRF_4_port, 
                           DATAIN(3) => MUXtoRF_3_port, DATAIN(2) => 
                           MUXtoRF_2_port, DATAIN(1) => MUXtoRF_1_port, 
                           DATAIN(0) => MUXtoRF_0_port, NPCfromIF(31) => 
                           NXPC_31_port, NPCfromIF(30) => NXPC_30_port, 
                           NPCfromIF(29) => NXPC_29_port, NPCfromIF(28) => 
                           NXPC_28_port, NPCfromIF(27) => NXPC_27_port, 
                           NPCfromIF(26) => NXPC_26_port, NPCfromIF(25) => 
                           NXPC_25_port, NPCfromIF(24) => NXPC_24_port, 
                           NPCfromIF(23) => NXPC_23_port, NPCfromIF(22) => 
                           NXPC_22_port, NPCfromIF(21) => NXPC_21_port, 
                           NPCfromIF(20) => NXPC_20_port, NPCfromIF(19) => 
                           NXPC_19_port, NPCfromIF(18) => NXPC_18_port, 
                           NPCfromIF(17) => NXPC_17_port, NPCfromIF(16) => 
                           NXPC_16_port, NPCfromIF(15) => NXPC_15_port, 
                           NPCfromIF(14) => NXPC_14_port, NPCfromIF(13) => 
                           NXPC_13_port, NPCfromIF(12) => NXPC_12_port, 
                           NPCfromIF(11) => NXPC_11_port, NPCfromIF(10) => 
                           NXPC_10_port, NPCfromIF(9) => NXPC_9_port, 
                           NPCfromIF(8) => NXPC_8_port, NPCfromIF(7) => 
                           NXPC_7_port, NPCfromIF(6) => NXPC_6_port, 
                           NPCfromIF(5) => NXPC_5_port, NPCfromIF(4) => 
                           NXPC_4_port, NPCfromIF(3) => NXPC_3_port, 
                           NPCfromIF(2) => NXPC_2_port, NPCfromIF(1) => 
                           NXPC_1_port, NPCfromIF(0) => NXPC_0_port, OUT1(31) 
                           => OUT1_31_port, OUT1(30) => OUT1_30_port, OUT1(29) 
                           => OUT1_29_port, OUT1(28) => OUT1_28_port, OUT1(27) 
                           => OUT1_27_port, OUT1(26) => OUT1_26_port, OUT1(25) 
                           => OUT1_25_port, OUT1(24) => OUT1_24_port, OUT1(23) 
                           => OUT1_23_port, OUT1(22) => OUT1_22_port, OUT1(21) 
                           => OUT1_21_port, OUT1(20) => OUT1_20_port, OUT1(19) 
                           => OUT1_19_port, OUT1(18) => OUT1_18_port, OUT1(17) 
                           => OUT1_17_port, OUT1(16) => OUT1_16_port, OUT1(15) 
                           => OUT1_15_port, OUT1(14) => OUT1_14_port, OUT1(13) 
                           => OUT1_13_port, OUT1(12) => OUT1_12_port, OUT1(11) 
                           => OUT1_11_port, OUT1(10) => OUT1_10_port, OUT1(9) 
                           => OUT1_9_port, OUT1(8) => OUT1_8_port, OUT1(7) => 
                           OUT1_7_port, OUT1(6) => OUT1_6_port, OUT1(5) => 
                           OUT1_5_port, OUT1(4) => OUT1_4_port, OUT1(3) => 
                           OUT1_3_port, OUT1(2) => OUT1_2_port, OUT1(1) => 
                           OUT1_1_port, OUT1(0) => OUT1_0_port, OUT2(31) => 
                           OUT2_31_port, OUT2(30) => OUT2_30_port, OUT2(29) => 
                           OUT2_29_port, OUT2(28) => OUT2_28_port, OUT2(27) => 
                           OUT2_27_port, OUT2(26) => OUT2_26_port, OUT2(25) => 
                           OUT2_25_port, OUT2(24) => OUT2_24_port, OUT2(23) => 
                           OUT2_23_port, OUT2(22) => OUT2_22_port, OUT2(21) => 
                           OUT2_21_port, OUT2(20) => OUT2_20_port, OUT2(19) => 
                           OUT2_19_port, OUT2(18) => OUT2_18_port, OUT2(17) => 
                           OUT2_17_port, OUT2(16) => OUT2_16_port, OUT2(15) => 
                           OUT2_15_port, OUT2(14) => OUT2_14_port, OUT2(13) => 
                           OUT2_13_port, OUT2(12) => OUT2_12_port, OUT2(11) => 
                           OUT2_11_port, OUT2(10) => OUT2_10_port, OUT2(9) => 
                           OUT2_9_port, OUT2(8) => OUT2_8_port, OUT2(7) => 
                           OUT2_7_port, OUT2(6) => OUT2_6_port, OUT2(5) => 
                           OUT2_5_port, OUT2(4) => OUT2_4_port, OUT2(3) => 
                           OUT2_3_port, OUT2(2) => OUT2_2_port, OUT2(1) => 
                           OUT2_1_port, OUT2(0) => OUT2_0_port, OUTNPC(31) => 
                           n_1354, OUTNPC(30) => n_1355, OUTNPC(29) => n_1356, 
                           OUTNPC(28) => n_1357, OUTNPC(27) => n_1358, 
                           OUTNPC(26) => n_1359, OUTNPC(25) => n_1360, 
                           OUTNPC(24) => n_1361, OUTNPC(23) => n_1362, 
                           OUTNPC(22) => n_1363, OUTNPC(21) => n_1364, 
                           OUTNPC(20) => n_1365, OUTNPC(19) => n_1366, 
                           OUTNPC(18) => n_1367, OUTNPC(17) => n_1368, 
                           OUTNPC(16) => n_1369, OUTNPC(15) => n_1370, 
                           OUTNPC(14) => n_1371, OUTNPC(13) => n_1372, 
                           OUTNPC(12) => n_1373, OUTNPC(11) => n_1374, 
                           OUTNPC(10) => n_1375, OUTNPC(9) => NewPC_9_port, 
                           OUTNPC(8) => NewPC_8_port, OUTNPC(7) => NewPC_7_port
                           , OUTNPC(6) => NewPC_6_port, OUTNPC(5) => 
                           NewPC_5_port, OUTNPC(4) => NewPC_4_port, OUTNPC(3) 
                           => NewPC_3_port, OUTNPC(2) => NewPC_2_port, 
                           OUTNPC(1) => NewPC_1_port, OUTNPC(0) => NewPC_0_port
                           , OUTIMM(31) => OUTIMM_31_port, OUTIMM(30) => 
                           OUTIMM_30_port, OUTIMM(29) => OUTIMM_29_port, 
                           OUTIMM(28) => OUTIMM_28_port, OUTIMM(27) => 
                           OUTIMM_27_port, OUTIMM(26) => OUTIMM_26_port, 
                           OUTIMM(25) => OUTIMM_25_port, OUTIMM(24) => 
                           OUTIMM_24_port, OUTIMM(23) => OUTIMM_23_port, 
                           OUTIMM(22) => OUTIMM_22_port, OUTIMM(21) => 
                           OUTIMM_21_port, OUTIMM(20) => OUTIMM_20_port, 
                           OUTIMM(19) => OUTIMM_19_port, OUTIMM(18) => 
                           OUTIMM_18_port, OUTIMM(17) => OUTIMM_17_port, 
                           OUTIMM(16) => OUTIMM_16_port, OUTIMM(15) => 
                           OUTIMM_15_port, OUTIMM(14) => OUTIMM_14_port, 
                           OUTIMM(13) => OUTIMM_13_port, OUTIMM(12) => 
                           OUTIMM_12_port, OUTIMM(11) => OUTIMM_11_port, 
                           OUTIMM(10) => OUTIMM_10_port, OUTIMM(9) => 
                           OUTIMM_9_port, OUTIMM(8) => OUTIMM_8_port, OUTIMM(7)
                           => OUTIMM_7_port, OUTIMM(6) => OUTIMM_6_port, 
                           OUTIMM(5) => OUTIMM_5_port, OUTIMM(4) => 
                           OUTIMM_4_port, OUTIMM(3) => OUTIMM_3_port, OUTIMM(2)
                           => OUTIMM_2_port, OUTIMM(1) => OUTIMM_1_port, 
                           OUTIMM(0) => OUTIMM_0_port, NPCtoEX(31) => 
                           NPCfromDECODE_31_port, NPCtoEX(30) => 
                           NPCfromDECODE_30_port, NPCtoEX(29) => 
                           NPCfromDECODE_29_port, NPCtoEX(28) => 
                           NPCfromDECODE_28_port, NPCtoEX(27) => 
                           NPCfromDECODE_27_port, NPCtoEX(26) => 
                           NPCfromDECODE_26_port, NPCtoEX(25) => 
                           NPCfromDECODE_25_port, NPCtoEX(24) => 
                           NPCfromDECODE_24_port, NPCtoEX(23) => 
                           NPCfromDECODE_23_port, NPCtoEX(22) => 
                           NPCfromDECODE_22_port, NPCtoEX(21) => 
                           NPCfromDECODE_21_port, NPCtoEX(20) => 
                           NPCfromDECODE_20_port, NPCtoEX(19) => 
                           NPCfromDECODE_19_port, NPCtoEX(18) => 
                           NPCfromDECODE_18_port, NPCtoEX(17) => 
                           NPCfromDECODE_17_port, NPCtoEX(16) => 
                           NPCfromDECODE_16_port, NPCtoEX(15) => 
                           NPCfromDECODE_15_port, NPCtoEX(14) => 
                           NPCfromDECODE_14_port, NPCtoEX(13) => 
                           NPCfromDECODE_13_port, NPCtoEX(12) => 
                           NPCfromDECODE_12_port, NPCtoEX(11) => 
                           NPCfromDECODE_11_port, NPCtoEX(10) => 
                           NPCfromDECODE_10_port, NPCtoEX(9) => 
                           NPCfromDECODE_9_port, NPCtoEX(8) => 
                           NPCfromDECODE_8_port, NPCtoEX(7) => 
                           NPCfromDECODE_7_port, NPCtoEX(6) => 
                           NPCfromDECODE_6_port, NPCtoEX(5) => 
                           NPCfromDECODE_5_port, NPCtoEX(4) => 
                           NPCfromDECODE_4_port, NPCtoEX(3) => 
                           NPCfromDECODE_3_port, NPCtoEX(2) => 
                           NPCfromDECODE_2_port, NPCtoEX(1) => 
                           NPCfromDECODE_1_port, NPCtoEX(0) => 
                           NPCfromDECODE_0_port, AddressWtoEX(31) => 
                           ADDWfromDECODE_31_port, AddressWtoEX(30) => 
                           ADDWfromDECODE_30_port, AddressWtoEX(29) => 
                           ADDWfromDECODE_29_port, AddressWtoEX(28) => 
                           ADDWfromDECODE_28_port, AddressWtoEX(27) => 
                           ADDWfromDECODE_27_port, AddressWtoEX(26) => 
                           ADDWfromDECODE_26_port, AddressWtoEX(25) => 
                           ADDWfromDECODE_25_port, AddressWtoEX(24) => 
                           ADDWfromDECODE_24_port, AddressWtoEX(23) => 
                           ADDWfromDECODE_23_port, AddressWtoEX(22) => 
                           ADDWfromDECODE_22_port, AddressWtoEX(21) => 
                           ADDWfromDECODE_21_port, AddressWtoEX(20) => 
                           ADDWfromDECODE_20_port, AddressWtoEX(19) => 
                           ADDWfromDECODE_19_port, AddressWtoEX(18) => 
                           ADDWfromDECODE_18_port, AddressWtoEX(17) => 
                           ADDWfromDECODE_17_port, AddressWtoEX(16) => 
                           ADDWfromDECODE_16_port, AddressWtoEX(15) => 
                           ADDWfromDECODE_15_port, AddressWtoEX(14) => 
                           ADDWfromDECODE_14_port, AddressWtoEX(13) => 
                           ADDWfromDECODE_13_port, AddressWtoEX(12) => 
                           ADDWfromDECODE_12_port, AddressWtoEX(11) => 
                           ADDWfromDECODE_11_port, AddressWtoEX(10) => 
                           ADDWfromDECODE_10_port, AddressWtoEX(9) => 
                           ADDWfromDECODE_9_port, AddressWtoEX(8) => 
                           ADDWfromDECODE_8_port, AddressWtoEX(7) => 
                           ADDWfromDECODE_7_port, AddressWtoEX(6) => 
                           ADDWfromDECODE_6_port, AddressWtoEX(5) => 
                           ADDWfromDECODE_5_port, AddressWtoEX(4) => 
                           ADDWfromDECODE_4_port, AddressWtoEX(3) => 
                           ADDWfromDECODE_3_port, AddressWtoEX(2) => 
                           ADDWfromDECODE_2_port, AddressWtoEX(1) => 
                           ADDWfromDECODE_1_port, AddressWtoEX(0) => 
                           ADDWfromDECODE_0_port, BRANCHtoFetch => 
                           BRANCHtoFetch);
   EU : executeUnit_M32_C4 port map( clock => clock, reset => n1, en3 => en3, 
                           Mux1Sel => Mux1Sel, Mux2Sel => Mux2Sel, ALUCODE(3) 
                           => ALUCODE(3), ALUCODE(2) => ALUCODE(2), ALUCODE(1) 
                           => ALUCODE(1), ALUCODE(0) => ALUCODE(0), OUT1RF(31) 
                           => OUT1_31_port, OUT1RF(30) => OUT1_30_port, 
                           OUT1RF(29) => OUT1_29_port, OUT1RF(28) => 
                           OUT1_28_port, OUT1RF(27) => OUT1_27_port, OUT1RF(26)
                           => OUT1_26_port, OUT1RF(25) => OUT1_25_port, 
                           OUT1RF(24) => OUT1_24_port, OUT1RF(23) => 
                           OUT1_23_port, OUT1RF(22) => OUT1_22_port, OUT1RF(21)
                           => OUT1_21_port, OUT1RF(20) => OUT1_20_port, 
                           OUT1RF(19) => OUT1_19_port, OUT1RF(18) => 
                           OUT1_18_port, OUT1RF(17) => OUT1_17_port, OUT1RF(16)
                           => OUT1_16_port, OUT1RF(15) => OUT1_15_port, 
                           OUT1RF(14) => OUT1_14_port, OUT1RF(13) => 
                           OUT1_13_port, OUT1RF(12) => OUT1_12_port, OUT1RF(11)
                           => OUT1_11_port, OUT1RF(10) => OUT1_10_port, 
                           OUT1RF(9) => OUT1_9_port, OUT1RF(8) => OUT1_8_port, 
                           OUT1RF(7) => OUT1_7_port, OUT1RF(6) => OUT1_6_port, 
                           OUT1RF(5) => OUT1_5_port, OUT1RF(4) => OUT1_4_port, 
                           OUT1RF(3) => OUT1_3_port, OUT1RF(2) => OUT1_2_port, 
                           OUT1RF(1) => OUT1_1_port, OUT1RF(0) => OUT1_0_port, 
                           OUT2RF(31) => OUT2_31_port, OUT2RF(30) => 
                           OUT2_30_port, OUT2RF(29) => OUT2_29_port, OUT2RF(28)
                           => OUT2_28_port, OUT2RF(27) => OUT2_27_port, 
                           OUT2RF(26) => OUT2_26_port, OUT2RF(25) => 
                           OUT2_25_port, OUT2RF(24) => OUT2_24_port, OUT2RF(23)
                           => OUT2_23_port, OUT2RF(22) => OUT2_22_port, 
                           OUT2RF(21) => OUT2_21_port, OUT2RF(20) => 
                           OUT2_20_port, OUT2RF(19) => OUT2_19_port, OUT2RF(18)
                           => OUT2_18_port, OUT2RF(17) => OUT2_17_port, 
                           OUT2RF(16) => OUT2_16_port, OUT2RF(15) => 
                           OUT2_15_port, OUT2RF(14) => OUT2_14_port, OUT2RF(13)
                           => OUT2_13_port, OUT2RF(12) => OUT2_12_port, 
                           OUT2RF(11) => OUT2_11_port, OUT2RF(10) => 
                           OUT2_10_port, OUT2RF(9) => OUT2_9_port, OUT2RF(8) =>
                           OUT2_8_port, OUT2RF(7) => OUT2_7_port, OUT2RF(6) => 
                           OUT2_6_port, OUT2RF(5) => OUT2_5_port, OUT2RF(4) => 
                           OUT2_4_port, OUT2RF(3) => OUT2_3_port, OUT2RF(2) => 
                           OUT2_2_port, OUT2RF(1) => OUT2_1_port, OUT2RF(0) => 
                           OUT2_0_port, IMMEDIATE(31) => OUTIMM_31_port, 
                           IMMEDIATE(30) => OUTIMM_30_port, IMMEDIATE(29) => 
                           OUTIMM_29_port, IMMEDIATE(28) => OUTIMM_28_port, 
                           IMMEDIATE(27) => OUTIMM_27_port, IMMEDIATE(26) => 
                           OUTIMM_26_port, IMMEDIATE(25) => OUTIMM_25_port, 
                           IMMEDIATE(24) => OUTIMM_24_port, IMMEDIATE(23) => 
                           OUTIMM_23_port, IMMEDIATE(22) => OUTIMM_22_port, 
                           IMMEDIATE(21) => OUTIMM_21_port, IMMEDIATE(20) => 
                           OUTIMM_20_port, IMMEDIATE(19) => OUTIMM_19_port, 
                           IMMEDIATE(18) => OUTIMM_18_port, IMMEDIATE(17) => 
                           OUTIMM_17_port, IMMEDIATE(16) => OUTIMM_16_port, 
                           IMMEDIATE(15) => OUTIMM_15_port, IMMEDIATE(14) => 
                           OUTIMM_14_port, IMMEDIATE(13) => OUTIMM_13_port, 
                           IMMEDIATE(12) => OUTIMM_12_port, IMMEDIATE(11) => 
                           OUTIMM_11_port, IMMEDIATE(10) => OUTIMM_10_port, 
                           IMMEDIATE(9) => OUTIMM_9_port, IMMEDIATE(8) => 
                           OUTIMM_8_port, IMMEDIATE(7) => OUTIMM_7_port, 
                           IMMEDIATE(6) => OUTIMM_6_port, IMMEDIATE(5) => 
                           OUTIMM_5_port, IMMEDIATE(4) => OUTIMM_4_port, 
                           IMMEDIATE(3) => OUTIMM_3_port, IMMEDIATE(2) => 
                           OUTIMM_2_port, IMMEDIATE(1) => OUTIMM_1_port, 
                           IMMEDIATE(0) => OUTIMM_0_port, NPCFromDecode(31) => 
                           NPCfromDECODE_31_port, NPCFromDecode(30) => 
                           NPCfromDECODE_30_port, NPCFromDecode(29) => 
                           NPCfromDECODE_29_port, NPCFromDecode(28) => 
                           NPCfromDECODE_28_port, NPCFromDecode(27) => 
                           NPCfromDECODE_27_port, NPCFromDecode(26) => 
                           NPCfromDECODE_26_port, NPCFromDecode(25) => 
                           NPCfromDECODE_25_port, NPCFromDecode(24) => 
                           NPCfromDECODE_24_port, NPCFromDecode(23) => 
                           NPCfromDECODE_23_port, NPCFromDecode(22) => 
                           NPCfromDECODE_22_port, NPCFromDecode(21) => 
                           NPCfromDECODE_21_port, NPCFromDecode(20) => 
                           NPCfromDECODE_20_port, NPCFromDecode(19) => 
                           NPCfromDECODE_19_port, NPCFromDecode(18) => 
                           NPCfromDECODE_18_port, NPCFromDecode(17) => 
                           NPCfromDECODE_17_port, NPCFromDecode(16) => 
                           NPCfromDECODE_16_port, NPCFromDecode(15) => 
                           NPCfromDECODE_15_port, NPCFromDecode(14) => 
                           NPCfromDECODE_14_port, NPCFromDecode(13) => 
                           NPCfromDECODE_13_port, NPCFromDecode(12) => 
                           NPCfromDECODE_12_port, NPCFromDecode(11) => 
                           NPCfromDECODE_11_port, NPCFromDecode(10) => 
                           NPCfromDECODE_10_port, NPCFromDecode(9) => 
                           NPCfromDECODE_9_port, NPCFromDecode(8) => 
                           NPCfromDECODE_8_port, NPCFromDecode(7) => 
                           NPCfromDECODE_7_port, NPCFromDecode(6) => 
                           NPCfromDECODE_6_port, NPCFromDecode(5) => 
                           NPCfromDECODE_5_port, NPCFromDecode(4) => 
                           NPCfromDECODE_4_port, NPCFromDecode(3) => 
                           NPCfromDECODE_3_port, NPCFromDecode(2) => 
                           NPCfromDECODE_2_port, NPCFromDecode(1) => 
                           NPCfromDECODE_1_port, NPCFromDecode(0) => 
                           NPCfromDECODE_0_port, AddressWfromDecode(31) => 
                           ADDWfromDECODE_31_port, AddressWfromDecode(30) => 
                           ADDWfromDECODE_30_port, AddressWfromDecode(29) => 
                           ADDWfromDECODE_29_port, AddressWfromDecode(28) => 
                           ADDWfromDECODE_28_port, AddressWfromDecode(27) => 
                           ADDWfromDECODE_27_port, AddressWfromDecode(26) => 
                           ADDWfromDECODE_26_port, AddressWfromDecode(25) => 
                           ADDWfromDECODE_25_port, AddressWfromDecode(24) => 
                           ADDWfromDECODE_24_port, AddressWfromDecode(23) => 
                           ADDWfromDECODE_23_port, AddressWfromDecode(22) => 
                           ADDWfromDECODE_22_port, AddressWfromDecode(21) => 
                           ADDWfromDECODE_21_port, AddressWfromDecode(20) => 
                           ADDWfromDECODE_20_port, AddressWfromDecode(19) => 
                           ADDWfromDECODE_19_port, AddressWfromDecode(18) => 
                           ADDWfromDECODE_18_port, AddressWfromDecode(17) => 
                           ADDWfromDECODE_17_port, AddressWfromDecode(16) => 
                           ADDWfromDECODE_16_port, AddressWfromDecode(15) => 
                           ADDWfromDECODE_15_port, AddressWfromDecode(14) => 
                           ADDWfromDECODE_14_port, AddressWfromDecode(13) => 
                           ADDWfromDECODE_13_port, AddressWfromDecode(12) => 
                           ADDWfromDECODE_12_port, AddressWfromDecode(11) => 
                           ADDWfromDECODE_11_port, AddressWfromDecode(10) => 
                           ADDWfromDECODE_10_port, AddressWfromDecode(9) => 
                           ADDWfromDECODE_9_port, AddressWfromDecode(8) => 
                           ADDWfromDECODE_8_port, AddressWfromDecode(7) => 
                           ADDWfromDECODE_7_port, AddressWfromDecode(6) => 
                           ADDWfromDECODE_6_port, AddressWfromDecode(5) => 
                           ADDWfromDECODE_5_port, AddressWfromDecode(4) => 
                           ADDWfromDECODE_4_port, AddressWfromDecode(3) => 
                           ADDWfromDECODE_3_port, AddressWfromDecode(2) => 
                           ADDWfromDECODE_2_port, AddressWfromDecode(1) => 
                           ADDWfromDECODE_1_port, AddressWfromDecode(0) => 
                           ADDWfromDECODE_0_port, ALUtoMEMORY(31) => 
                           ALUtoMEMORY_31_port, ALUtoMEMORY(30) => 
                           ALUtoMEMORY_30_port, ALUtoMEMORY(29) => 
                           ALUtoMEMORY_29_port, ALUtoMEMORY(28) => 
                           ALUtoMEMORY_28_port, ALUtoMEMORY(27) => 
                           ALUtoMEMORY_27_port, ALUtoMEMORY(26) => 
                           ALUtoMEMORY_26_port, ALUtoMEMORY(25) => 
                           ALUtoMEMORY_25_port, ALUtoMEMORY(24) => 
                           ALUtoMEMORY_24_port, ALUtoMEMORY(23) => 
                           ALUtoMEMORY_23_port, ALUtoMEMORY(22) => 
                           ALUtoMEMORY_22_port, ALUtoMEMORY(21) => 
                           ALUtoMEMORY_21_port, ALUtoMEMORY(20) => 
                           ALUtoMEMORY_20_port, ALUtoMEMORY(19) => 
                           ALUtoMEMORY_19_port, ALUtoMEMORY(18) => 
                           ALUtoMEMORY_18_port, ALUtoMEMORY(17) => 
                           ALUtoMEMORY_17_port, ALUtoMEMORY(16) => 
                           ALUtoMEMORY_16_port, ALUtoMEMORY(15) => 
                           ALUtoMEMORY_15_port, ALUtoMEMORY(14) => 
                           ALUtoMEMORY_14_port, ALUtoMEMORY(13) => 
                           ALUtoMEMORY_13_port, ALUtoMEMORY(12) => 
                           ALUtoMEMORY_12_port, ALUtoMEMORY(11) => 
                           ALUtoMEMORY_11_port, ALUtoMEMORY(10) => 
                           ALUtoMEMORY_10_port, ALUtoMEMORY(9) => 
                           ALUtoMEMORY_9_port, ALUtoMEMORY(8) => 
                           ALUtoMEMORY_8_port, ALUtoMEMORY(7) => 
                           ALUtoMEMORY_7_port, ALUtoMEMORY(6) => 
                           ALUtoMEMORY_6_port, ALUtoMEMORY(5) => 
                           ALUtoMEMORY_5_port, ALUtoMEMORY(4) => 
                           ALUtoMEMORY_4_port, ALUtoMEMORY(3) => 
                           ALUtoMEMORY_3_port, ALUtoMEMORY(2) => 
                           ALUtoMEMORY_2_port, ALUtoMEMORY(1) => 
                           ALUtoMEMORY_1_port, ALUtoMEMORY(0) => 
                           ALUtoMEMORY_0_port, OUT2RFtoMEMORY(31) => 
                           OUT2RFtoMEMORY(31), OUT2RFtoMEMORY(30) => 
                           OUT2RFtoMEMORY(30), OUT2RFtoMEMORY(29) => 
                           OUT2RFtoMEMORY(29), OUT2RFtoMEMORY(28) => 
                           OUT2RFtoMEMORY(28), OUT2RFtoMEMORY(27) => 
                           OUT2RFtoMEMORY(27), OUT2RFtoMEMORY(26) => 
                           OUT2RFtoMEMORY(26), OUT2RFtoMEMORY(25) => 
                           OUT2RFtoMEMORY(25), OUT2RFtoMEMORY(24) => 
                           OUT2RFtoMEMORY(24), OUT2RFtoMEMORY(23) => 
                           OUT2RFtoMEMORY(23), OUT2RFtoMEMORY(22) => 
                           OUT2RFtoMEMORY(22), OUT2RFtoMEMORY(21) => 
                           OUT2RFtoMEMORY(21), OUT2RFtoMEMORY(20) => 
                           OUT2RFtoMEMORY(20), OUT2RFtoMEMORY(19) => 
                           OUT2RFtoMEMORY(19), OUT2RFtoMEMORY(18) => 
                           OUT2RFtoMEMORY(18), OUT2RFtoMEMORY(17) => 
                           OUT2RFtoMEMORY(17), OUT2RFtoMEMORY(16) => 
                           OUT2RFtoMEMORY(16), OUT2RFtoMEMORY(15) => 
                           OUT2RFtoMEMORY(15), OUT2RFtoMEMORY(14) => 
                           OUT2RFtoMEMORY(14), OUT2RFtoMEMORY(13) => 
                           OUT2RFtoMEMORY(13), OUT2RFtoMEMORY(12) => 
                           OUT2RFtoMEMORY(12), OUT2RFtoMEMORY(11) => 
                           OUT2RFtoMEMORY(11), OUT2RFtoMEMORY(10) => 
                           OUT2RFtoMEMORY(10), OUT2RFtoMEMORY(9) => 
                           OUT2RFtoMEMORY(9), OUT2RFtoMEMORY(8) => 
                           OUT2RFtoMEMORY(8), OUT2RFtoMEMORY(7) => 
                           OUT2RFtoMEMORY(7), OUT2RFtoMEMORY(6) => 
                           OUT2RFtoMEMORY(6), OUT2RFtoMEMORY(5) => 
                           OUT2RFtoMEMORY(5), OUT2RFtoMEMORY(4) => 
                           OUT2RFtoMEMORY(4), OUT2RFtoMEMORY(3) => 
                           OUT2RFtoMEMORY(3), OUT2RFtoMEMORY(2) => 
                           OUT2RFtoMEMORY(2), OUT2RFtoMEMORY(1) => 
                           OUT2RFtoMEMORY(1), OUT2RFtoMEMORY(0) => 
                           OUT2RFtoMEMORY(0), AddressWtoMEMORY(31) => 
                           ADDWtoMEMORY_31_port, AddressWtoMEMORY(30) => 
                           ADDWtoMEMORY_30_port, AddressWtoMEMORY(29) => 
                           ADDWtoMEMORY_29_port, AddressWtoMEMORY(28) => 
                           ADDWtoMEMORY_28_port, AddressWtoMEMORY(27) => 
                           ADDWtoMEMORY_27_port, AddressWtoMEMORY(26) => 
                           ADDWtoMEMORY_26_port, AddressWtoMEMORY(25) => 
                           ADDWtoMEMORY_25_port, AddressWtoMEMORY(24) => 
                           ADDWtoMEMORY_24_port, AddressWtoMEMORY(23) => 
                           ADDWtoMEMORY_23_port, AddressWtoMEMORY(22) => 
                           ADDWtoMEMORY_22_port, AddressWtoMEMORY(21) => 
                           ADDWtoMEMORY_21_port, AddressWtoMEMORY(20) => 
                           ADDWtoMEMORY_20_port, AddressWtoMEMORY(19) => 
                           ADDWtoMEMORY_19_port, AddressWtoMEMORY(18) => 
                           ADDWtoMEMORY_18_port, AddressWtoMEMORY(17) => 
                           ADDWtoMEMORY_17_port, AddressWtoMEMORY(16) => 
                           ADDWtoMEMORY_16_port, AddressWtoMEMORY(15) => 
                           ADDWtoMEMORY_15_port, AddressWtoMEMORY(14) => 
                           ADDWtoMEMORY_14_port, AddressWtoMEMORY(13) => 
                           ADDWtoMEMORY_13_port, AddressWtoMEMORY(12) => 
                           ADDWtoMEMORY_12_port, AddressWtoMEMORY(11) => 
                           ADDWtoMEMORY_11_port, AddressWtoMEMORY(10) => 
                           ADDWtoMEMORY_10_port, AddressWtoMEMORY(9) => 
                           ADDWtoMEMORY_9_port, AddressWtoMEMORY(8) => 
                           ADDWtoMEMORY_8_port, AddressWtoMEMORY(7) => 
                           ADDWtoMEMORY_7_port, AddressWtoMEMORY(6) => 
                           ADDWtoMEMORY_6_port, AddressWtoMEMORY(5) => 
                           ADDWtoMEMORY_5_port, AddressWtoMEMORY(4) => 
                           ADDWtoMEMORY_4_port, AddressWtoMEMORY(3) => 
                           ADDWtoMEMORY_3_port, AddressWtoMEMORY(2) => 
                           ADDWtoMEMORY_2_port, AddressWtoMEMORY(1) => 
                           ADDWtoMEMORY_1_port, AddressWtoMEMORY(0) => 
                           ADDWtoMEMORY_0_port);
   MU : memoryUnit port map( clock => clock, reset => n1, en4 => en4, 
                           ALUout(31) => ALUtoMEMORY_31_port, ALUout(30) => 
                           ALUtoMEMORY_30_port, ALUout(29) => 
                           ALUtoMEMORY_29_port, ALUout(28) => 
                           ALUtoMEMORY_28_port, ALUout(27) => 
                           ALUtoMEMORY_27_port, ALUout(26) => 
                           ALUtoMEMORY_26_port, ALUout(25) => 
                           ALUtoMEMORY_25_port, ALUout(24) => 
                           ALUtoMEMORY_24_port, ALUout(23) => 
                           ALUtoMEMORY_23_port, ALUout(22) => 
                           ALUtoMEMORY_22_port, ALUout(21) => 
                           ALUtoMEMORY_21_port, ALUout(20) => 
                           ALUtoMEMORY_20_port, ALUout(19) => 
                           ALUtoMEMORY_19_port, ALUout(18) => 
                           ALUtoMEMORY_18_port, ALUout(17) => 
                           ALUtoMEMORY_17_port, ALUout(16) => 
                           ALUtoMEMORY_16_port, ALUout(15) => 
                           ALUtoMEMORY_15_port, ALUout(14) => 
                           ALUtoMEMORY_14_port, ALUout(13) => 
                           ALUtoMEMORY_13_port, ALUout(12) => 
                           ALUtoMEMORY_12_port, ALUout(11) => 
                           ALUtoMEMORY_11_port, ALUout(10) => 
                           ALUtoMEMORY_10_port, ALUout(9) => ALUtoMEMORY_9_port
                           , ALUout(8) => ALUtoMEMORY_8_port, ALUout(7) => 
                           ALUtoMEMORY_7_port, ALUout(6) => ALUtoMEMORY_6_port,
                           ALUout(5) => ALUtoMEMORY_5_port, ALUout(4) => 
                           ALUtoMEMORY_4_port, ALUout(3) => ALUtoMEMORY_3_port,
                           ALUout(2) => ALUtoMEMORY_2_port, ALUout(1) => 
                           ALUtoMEMORY_1_port, ALUout(0) => ALUtoMEMORY_0_port,
                           DRAMout(31) => DRAMout(31), DRAMout(30) => 
                           DRAMout(30), DRAMout(29) => DRAMout(29), DRAMout(28)
                           => DRAMout(28), DRAMout(27) => DRAMout(27), 
                           DRAMout(26) => DRAMout(26), DRAMout(25) => 
                           DRAMout(25), DRAMout(24) => DRAMout(24), DRAMout(23)
                           => DRAMout(23), DRAMout(22) => DRAMout(22), 
                           DRAMout(21) => DRAMout(21), DRAMout(20) => 
                           DRAMout(20), DRAMout(19) => DRAMout(19), DRAMout(18)
                           => DRAMout(18), DRAMout(17) => DRAMout(17), 
                           DRAMout(16) => DRAMout(16), DRAMout(15) => 
                           DRAMout(15), DRAMout(14) => DRAMout(14), DRAMout(13)
                           => DRAMout(13), DRAMout(12) => DRAMout(12), 
                           DRAMout(11) => DRAMout(11), DRAMout(10) => 
                           DRAMout(10), DRAMout(9) => DRAMout(9), DRAMout(8) =>
                           DRAMout(8), DRAMout(7) => DRAMout(7), DRAMout(6) => 
                           DRAMout(6), DRAMout(5) => DRAMout(5), DRAMout(4) => 
                           DRAMout(4), DRAMout(3) => DRAMout(3), DRAMout(2) => 
                           DRAMout(2), DRAMout(1) => DRAMout(1), DRAMout(0) => 
                           DRAMout(0), AddressWfromEXECUTE(31) => 
                           ADDWtoMEMORY_31_port, AddressWfromEXECUTE(30) => 
                           ADDWtoMEMORY_30_port, AddressWfromEXECUTE(29) => 
                           ADDWtoMEMORY_29_port, AddressWfromEXECUTE(28) => 
                           ADDWtoMEMORY_28_port, AddressWfromEXECUTE(27) => 
                           ADDWtoMEMORY_27_port, AddressWfromEXECUTE(26) => 
                           ADDWtoMEMORY_26_port, AddressWfromEXECUTE(25) => 
                           ADDWtoMEMORY_25_port, AddressWfromEXECUTE(24) => 
                           ADDWtoMEMORY_24_port, AddressWfromEXECUTE(23) => 
                           ADDWtoMEMORY_23_port, AddressWfromEXECUTE(22) => 
                           ADDWtoMEMORY_22_port, AddressWfromEXECUTE(21) => 
                           ADDWtoMEMORY_21_port, AddressWfromEXECUTE(20) => 
                           ADDWtoMEMORY_20_port, AddressWfromEXECUTE(19) => 
                           ADDWtoMEMORY_19_port, AddressWfromEXECUTE(18) => 
                           ADDWtoMEMORY_18_port, AddressWfromEXECUTE(17) => 
                           ADDWtoMEMORY_17_port, AddressWfromEXECUTE(16) => 
                           ADDWtoMEMORY_16_port, AddressWfromEXECUTE(15) => 
                           ADDWtoMEMORY_15_port, AddressWfromEXECUTE(14) => 
                           ADDWtoMEMORY_14_port, AddressWfromEXECUTE(13) => 
                           ADDWtoMEMORY_13_port, AddressWfromEXECUTE(12) => 
                           ADDWtoMEMORY_12_port, AddressWfromEXECUTE(11) => 
                           ADDWtoMEMORY_11_port, AddressWfromEXECUTE(10) => 
                           ADDWtoMEMORY_10_port, AddressWfromEXECUTE(9) => 
                           ADDWtoMEMORY_9_port, AddressWfromEXECUTE(8) => 
                           ADDWtoMEMORY_8_port, AddressWfromEXECUTE(7) => 
                           ADDWtoMEMORY_7_port, AddressWfromEXECUTE(6) => 
                           ADDWtoMEMORY_6_port, AddressWfromEXECUTE(5) => 
                           ADDWtoMEMORY_5_port, AddressWfromEXECUTE(4) => 
                           ADDWtoMEMORY_4_port, AddressWfromEXECUTE(3) => 
                           ADDWtoMEMORY_3_port, AddressWfromEXECUTE(2) => 
                           ADDWtoMEMORY_2_port, AddressWfromEXECUTE(1) => 
                           ADDWtoMEMORY_1_port, AddressWfromEXECUTE(0) => 
                           ADDWtoMEMORY_0_port, LOADDATA(31) => 
                           LOADDATA_31_port, LOADDATA(30) => LOADDATA_30_port, 
                           LOADDATA(29) => LOADDATA_29_port, LOADDATA(28) => 
                           LOADDATA_28_port, LOADDATA(27) => LOADDATA_27_port, 
                           LOADDATA(26) => LOADDATA_26_port, LOADDATA(25) => 
                           LOADDATA_25_port, LOADDATA(24) => LOADDATA_24_port, 
                           LOADDATA(23) => LOADDATA_23_port, LOADDATA(22) => 
                           LOADDATA_22_port, LOADDATA(21) => LOADDATA_21_port, 
                           LOADDATA(20) => LOADDATA_20_port, LOADDATA(19) => 
                           LOADDATA_19_port, LOADDATA(18) => LOADDATA_18_port, 
                           LOADDATA(17) => LOADDATA_17_port, LOADDATA(16) => 
                           LOADDATA_16_port, LOADDATA(15) => LOADDATA_15_port, 
                           LOADDATA(14) => LOADDATA_14_port, LOADDATA(13) => 
                           LOADDATA_13_port, LOADDATA(12) => LOADDATA_12_port, 
                           LOADDATA(11) => LOADDATA_11_port, LOADDATA(10) => 
                           LOADDATA_10_port, LOADDATA(9) => LOADDATA_9_port, 
                           LOADDATA(8) => LOADDATA_8_port, LOADDATA(7) => 
                           LOADDATA_7_port, LOADDATA(6) => LOADDATA_6_port, 
                           LOADDATA(5) => LOADDATA_5_port, LOADDATA(4) => 
                           LOADDATA_4_port, LOADDATA(3) => LOADDATA_3_port, 
                           LOADDATA(2) => LOADDATA_2_port, LOADDATA(1) => 
                           LOADDATA_1_port, LOADDATA(0) => LOADDATA_0_port, 
                           ALUtoWBMUX(31) => ALUtoWBMUX_31_port, ALUtoWBMUX(30)
                           => ALUtoWBMUX_30_port, ALUtoWBMUX(29) => 
                           ALUtoWBMUX_29_port, ALUtoWBMUX(28) => 
                           ALUtoWBMUX_28_port, ALUtoWBMUX(27) => 
                           ALUtoWBMUX_27_port, ALUtoWBMUX(26) => 
                           ALUtoWBMUX_26_port, ALUtoWBMUX(25) => 
                           ALUtoWBMUX_25_port, ALUtoWBMUX(24) => 
                           ALUtoWBMUX_24_port, ALUtoWBMUX(23) => 
                           ALUtoWBMUX_23_port, ALUtoWBMUX(22) => 
                           ALUtoWBMUX_22_port, ALUtoWBMUX(21) => 
                           ALUtoWBMUX_21_port, ALUtoWBMUX(20) => 
                           ALUtoWBMUX_20_port, ALUtoWBMUX(19) => 
                           ALUtoWBMUX_19_port, ALUtoWBMUX(18) => 
                           ALUtoWBMUX_18_port, ALUtoWBMUX(17) => 
                           ALUtoWBMUX_17_port, ALUtoWBMUX(16) => 
                           ALUtoWBMUX_16_port, ALUtoWBMUX(15) => 
                           ALUtoWBMUX_15_port, ALUtoWBMUX(14) => 
                           ALUtoWBMUX_14_port, ALUtoWBMUX(13) => 
                           ALUtoWBMUX_13_port, ALUtoWBMUX(12) => 
                           ALUtoWBMUX_12_port, ALUtoWBMUX(11) => 
                           ALUtoWBMUX_11_port, ALUtoWBMUX(10) => 
                           ALUtoWBMUX_10_port, ALUtoWBMUX(9) => 
                           ALUtoWBMUX_9_port, ALUtoWBMUX(8) => 
                           ALUtoWBMUX_8_port, ALUtoWBMUX(7) => 
                           ALUtoWBMUX_7_port, ALUtoWBMUX(6) => 
                           ALUtoWBMUX_6_port, ALUtoWBMUX(5) => 
                           ALUtoWBMUX_5_port, ALUtoWBMUX(4) => 
                           ALUtoWBMUX_4_port, ALUtoWBMUX(3) => 
                           ALUtoWBMUX_3_port, ALUtoWBMUX(2) => 
                           ALUtoWBMUX_2_port, ALUtoWBMUX(1) => 
                           ALUtoWBMUX_1_port, ALUtoWBMUX(0) => 
                           ALUtoWBMUX_0_port, AddressWtoWB(31) => 
                           ADDWtoWB_31_port, AddressWtoWB(30) => 
                           ADDWtoWB_30_port, AddressWtoWB(29) => 
                           ADDWtoWB_29_port, AddressWtoWB(28) => 
                           ADDWtoWB_28_port, AddressWtoWB(27) => 
                           ADDWtoWB_27_port, AddressWtoWB(26) => 
                           ADDWtoWB_26_port, AddressWtoWB(25) => 
                           ADDWtoWB_25_port, AddressWtoWB(24) => 
                           ADDWtoWB_24_port, AddressWtoWB(23) => 
                           ADDWtoWB_23_port, AddressWtoWB(22) => 
                           ADDWtoWB_22_port, AddressWtoWB(21) => 
                           ADDWtoWB_21_port, AddressWtoWB(20) => 
                           ADDWtoWB_20_port, AddressWtoWB(19) => 
                           ADDWtoWB_19_port, AddressWtoWB(18) => 
                           ADDWtoWB_18_port, AddressWtoWB(17) => 
                           ADDWtoWB_17_port, AddressWtoWB(16) => 
                           ADDWtoWB_16_port, AddressWtoWB(15) => 
                           ADDWtoWB_15_port, AddressWtoWB(14) => 
                           ADDWtoWB_14_port, AddressWtoWB(13) => 
                           ADDWtoWB_13_port, AddressWtoWB(12) => 
                           ADDWtoWB_12_port, AddressWtoWB(11) => 
                           ADDWtoWB_11_port, AddressWtoWB(10) => 
                           ADDWtoWB_10_port, AddressWtoWB(9) => ADDWtoWB_9_port
                           , AddressWtoWB(8) => ADDWtoWB_8_port, 
                           AddressWtoWB(7) => ADDWtoWB_7_port, AddressWtoWB(6) 
                           => ADDWtoWB_6_port, AddressWtoWB(5) => 
                           ADDWtoWB_5_port, AddressWtoWB(4) => ADDWtoWB_4_port,
                           AddressWtoWB(3) => ADDWtoWB_3_port, AddressWtoWB(2) 
                           => ADDWtoWB_2_port, AddressWtoWB(1) => 
                           ADDWtoWB_1_port, AddressWtoWB(0) => ADDWtoWB_0_port)
                           ;
   WBU : WBUnit port map( selwb => selwb, ALUin(31) => ALUtoWBMUX_31_port, 
                           ALUin(30) => ALUtoWBMUX_30_port, ALUin(29) => 
                           ALUtoWBMUX_29_port, ALUin(28) => ALUtoWBMUX_28_port,
                           ALUin(27) => ALUtoWBMUX_27_port, ALUin(26) => 
                           ALUtoWBMUX_26_port, ALUin(25) => ALUtoWBMUX_25_port,
                           ALUin(24) => ALUtoWBMUX_24_port, ALUin(23) => 
                           ALUtoWBMUX_23_port, ALUin(22) => ALUtoWBMUX_22_port,
                           ALUin(21) => ALUtoWBMUX_21_port, ALUin(20) => 
                           ALUtoWBMUX_20_port, ALUin(19) => ALUtoWBMUX_19_port,
                           ALUin(18) => ALUtoWBMUX_18_port, ALUin(17) => 
                           ALUtoWBMUX_17_port, ALUin(16) => ALUtoWBMUX_16_port,
                           ALUin(15) => ALUtoWBMUX_15_port, ALUin(14) => 
                           ALUtoWBMUX_14_port, ALUin(13) => ALUtoWBMUX_13_port,
                           ALUin(12) => ALUtoWBMUX_12_port, ALUin(11) => 
                           ALUtoWBMUX_11_port, ALUin(10) => ALUtoWBMUX_10_port,
                           ALUin(9) => ALUtoWBMUX_9_port, ALUin(8) => 
                           ALUtoWBMUX_8_port, ALUin(7) => ALUtoWBMUX_7_port, 
                           ALUin(6) => ALUtoWBMUX_6_port, ALUin(5) => 
                           ALUtoWBMUX_5_port, ALUin(4) => ALUtoWBMUX_4_port, 
                           ALUin(3) => ALUtoWBMUX_3_port, ALUin(2) => 
                           ALUtoWBMUX_2_port, ALUin(1) => ALUtoWBMUX_1_port, 
                           ALUin(0) => ALUtoWBMUX_0_port, LOADDATA(31) => 
                           LOADDATA_31_port, LOADDATA(30) => LOADDATA_30_port, 
                           LOADDATA(29) => LOADDATA_29_port, LOADDATA(28) => 
                           LOADDATA_28_port, LOADDATA(27) => LOADDATA_27_port, 
                           LOADDATA(26) => LOADDATA_26_port, LOADDATA(25) => 
                           LOADDATA_25_port, LOADDATA(24) => LOADDATA_24_port, 
                           LOADDATA(23) => LOADDATA_23_port, LOADDATA(22) => 
                           LOADDATA_22_port, LOADDATA(21) => LOADDATA_21_port, 
                           LOADDATA(20) => LOADDATA_20_port, LOADDATA(19) => 
                           LOADDATA_19_port, LOADDATA(18) => LOADDATA_18_port, 
                           LOADDATA(17) => LOADDATA_17_port, LOADDATA(16) => 
                           LOADDATA_16_port, LOADDATA(15) => LOADDATA_15_port, 
                           LOADDATA(14) => LOADDATA_14_port, LOADDATA(13) => 
                           LOADDATA_13_port, LOADDATA(12) => LOADDATA_12_port, 
                           LOADDATA(11) => LOADDATA_11_port, LOADDATA(10) => 
                           LOADDATA_10_port, LOADDATA(9) => LOADDATA_9_port, 
                           LOADDATA(8) => LOADDATA_8_port, LOADDATA(7) => 
                           LOADDATA_7_port, LOADDATA(6) => LOADDATA_6_port, 
                           LOADDATA(5) => LOADDATA_5_port, LOADDATA(4) => 
                           LOADDATA_4_port, LOADDATA(3) => LOADDATA_3_port, 
                           LOADDATA(2) => LOADDATA_2_port, LOADDATA(1) => 
                           LOADDATA_1_port, LOADDATA(0) => LOADDATA_0_port, 
                           AddressWfromMemory(31) => ADDWtoWB_31_port, 
                           AddressWfromMemory(30) => ADDWtoWB_30_port, 
                           AddressWfromMemory(29) => ADDWtoWB_29_port, 
                           AddressWfromMemory(28) => ADDWtoWB_28_port, 
                           AddressWfromMemory(27) => ADDWtoWB_27_port, 
                           AddressWfromMemory(26) => ADDWtoWB_26_port, 
                           AddressWfromMemory(25) => ADDWtoWB_25_port, 
                           AddressWfromMemory(24) => ADDWtoWB_24_port, 
                           AddressWfromMemory(23) => ADDWtoWB_23_port, 
                           AddressWfromMemory(22) => ADDWtoWB_22_port, 
                           AddressWfromMemory(21) => ADDWtoWB_21_port, 
                           AddressWfromMemory(20) => ADDWtoWB_20_port, 
                           AddressWfromMemory(19) => ADDWtoWB_19_port, 
                           AddressWfromMemory(18) => ADDWtoWB_18_port, 
                           AddressWfromMemory(17) => ADDWtoWB_17_port, 
                           AddressWfromMemory(16) => ADDWtoWB_16_port, 
                           AddressWfromMemory(15) => ADDWtoWB_15_port, 
                           AddressWfromMemory(14) => ADDWtoWB_14_port, 
                           AddressWfromMemory(13) => ADDWtoWB_13_port, 
                           AddressWfromMemory(12) => ADDWtoWB_12_port, 
                           AddressWfromMemory(11) => ADDWtoWB_11_port, 
                           AddressWfromMemory(10) => ADDWtoWB_10_port, 
                           AddressWfromMemory(9) => ADDWtoWB_9_port, 
                           AddressWfromMemory(8) => ADDWtoWB_8_port, 
                           AddressWfromMemory(7) => ADDWtoWB_7_port, 
                           AddressWfromMemory(6) => ADDWtoWB_6_port, 
                           AddressWfromMemory(5) => ADDWtoWB_5_port, 
                           AddressWfromMemory(4) => ADDWtoWB_4_port, 
                           AddressWfromMemory(3) => ADDWtoWB_3_port, 
                           AddressWfromMemory(2) => ADDWtoWB_2_port, 
                           AddressWfromMemory(1) => ADDWtoWB_1_port, 
                           AddressWfromMemory(0) => ADDWtoWB_0_port, 
                           MUXtoRF(31) => MUXtoRF_31_port, MUXtoRF(30) => 
                           MUXtoRF_30_port, MUXtoRF(29) => MUXtoRF_29_port, 
                           MUXtoRF(28) => MUXtoRF_28_port, MUXtoRF(27) => 
                           MUXtoRF_27_port, MUXtoRF(26) => MUXtoRF_26_port, 
                           MUXtoRF(25) => MUXtoRF_25_port, MUXtoRF(24) => 
                           MUXtoRF_24_port, MUXtoRF(23) => MUXtoRF_23_port, 
                           MUXtoRF(22) => MUXtoRF_22_port, MUXtoRF(21) => 
                           MUXtoRF_21_port, MUXtoRF(20) => MUXtoRF_20_port, 
                           MUXtoRF(19) => MUXtoRF_19_port, MUXtoRF(18) => 
                           MUXtoRF_18_port, MUXtoRF(17) => MUXtoRF_17_port, 
                           MUXtoRF(16) => MUXtoRF_16_port, MUXtoRF(15) => 
                           MUXtoRF_15_port, MUXtoRF(14) => MUXtoRF_14_port, 
                           MUXtoRF(13) => MUXtoRF_13_port, MUXtoRF(12) => 
                           MUXtoRF_12_port, MUXtoRF(11) => MUXtoRF_11_port, 
                           MUXtoRF(10) => MUXtoRF_10_port, MUXtoRF(9) => 
                           MUXtoRF_9_port, MUXtoRF(8) => MUXtoRF_8_port, 
                           MUXtoRF(7) => MUXtoRF_7_port, MUXtoRF(6) => 
                           MUXtoRF_6_port, MUXtoRF(5) => MUXtoRF_5_port, 
                           MUXtoRF(4) => MUXtoRF_4_port, MUXtoRF(3) => 
                           MUXtoRF_3_port, MUXtoRF(2) => MUXtoRF_2_port, 
                           MUXtoRF(1) => MUXtoRF_1_port, MUXtoRF(0) => 
                           MUXtoRF_0_port, AddressWtoDECODE(31) => n_1376, 
                           AddressWtoDECODE(30) => n_1377, AddressWtoDECODE(29)
                           => n_1378, AddressWtoDECODE(28) => n_1379, 
                           AddressWtoDECODE(27) => n_1380, AddressWtoDECODE(26)
                           => n_1381, AddressWtoDECODE(25) => n_1382, 
                           AddressWtoDECODE(24) => n_1383, AddressWtoDECODE(23)
                           => n_1384, AddressWtoDECODE(22) => n_1385, 
                           AddressWtoDECODE(21) => n_1386, AddressWtoDECODE(20)
                           => n_1387, AddressWtoDECODE(19) => n_1388, 
                           AddressWtoDECODE(18) => n_1389, AddressWtoDECODE(17)
                           => n_1390, AddressWtoDECODE(16) => n_1391, 
                           AddressWtoDECODE(15) => n_1392, AddressWtoDECODE(14)
                           => n_1393, AddressWtoDECODE(13) => n_1394, 
                           AddressWtoDECODE(12) => n_1395, AddressWtoDECODE(11)
                           => n_1396, AddressWtoDECODE(10) => n_1397, 
                           AddressWtoDECODE(9) => n_1398, AddressWtoDECODE(8) 
                           => n_1399, AddressWtoDECODE(7) => n_1400, 
                           AddressWtoDECODE(6) => n_1401, AddressWtoDECODE(5) 
                           => n_1402, AddressWtoDECODE(4) => 
                           AddressfromWB_4_port, AddressWtoDECODE(3) => 
                           AddressfromWB_3_port, AddressWtoDECODE(2) => 
                           AddressfromWB_2_port, AddressWtoDECODE(1) => 
                           AddressfromWB_1_port, AddressWtoDECODE(0) => 
                           AddressfromWB_0_port);
   U23 : BUF_X1 port map( A => reset, Z => n1);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         en1, en2, SignSelect, RD1, RD2, JMP, BranchCondSel, BRANCHenable, 
         RegDestination, en3, Mux1Sel, Mux2Sel : out std_logic;  ALUCODE : out 
         std_logic_vector (3 downto 0);  en4, MemoryEnable, ReadNotWrite, selwb
         , WR : out std_logic);

end Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17;

architecture SYN_structural of 
   Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal ALUCODE_3_port, ALUCODE_2_port, ALUCODE_1_port, ALUCODE_0_port, 
      cw2_7_port, cw2_6_port, cw2_5_port, cw2_4_port, cw2_3_port, cw2_2_port, 
      cw2_1_port, cw2_0_port, N174, N175, N176, N182, N183, N184, N185, n3, n6,
      n8, n10, n12, n13, n14, n15, n103, n104, n105, n193, n194, n195, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n358, n359, n360, n361, 
      n362, n364, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n363, n365, n366, n367, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
      n95, n96, n97, n98, n99, n100, n101, n102, n106, n107, n108, n109, n110, 
      n111, n112, n113, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409,
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418 : 
      std_logic;

begin
   ALUCODE <= ( ALUCODE_3_port, ALUCODE_2_port, ALUCODE_1_port, ALUCODE_0_port 
      );
   
   en1 <= '1';
   aluOpcode3_reg_3_inst : DFF_X1 port map( D => n105, CK => Clk, Q => 
                           ALUCODE_3_port, QN => n195);
   aluOpcode3_reg_2_inst : DFF_X1 port map( D => n104, CK => Clk, Q => 
                           ALUCODE_2_port, QN => n194);
   aluOpcode3_reg_1_inst : DFF_X1 port map( D => n87, CK => Clk, Q => 
                           ALUCODE_1_port, QN => n_1403);
   cw2_reg_15_inst : DLH_X1 port map( G => N174, D => n85, Q => en2);
   cw2_reg_13_inst : DLH_X1 port map( G => N174, D => N184, Q => RD1);
   cw2_reg_12_inst : DLH_X1 port map( G => N174, D => N183, Q => RD2);
   cw2_reg_11_inst : DLH_X1 port map( G => N174, D => N182, Q => JMP);
   cw2_reg_10_inst : DLH_X1 port map( G => N174, D => n364, Q => BranchCondSel)
                           ;
   cw2_reg_9_inst : DLH_X1 port map( G => N174, D => n90, Q => BRANCHenable);
   cw2_reg_8_inst : DLH_X1 port map( G => N174, D => n88, Q => RegDestination);
   cw2_reg_7_inst : DLH_X1 port map( G => N174, D => n85, Q => cw2_7_port);
   cw3_reg_7_inst : SDFF_X1 port map( D => n15, SI => n85, SE => cw2_7_port, CK
                           => Clk, Q => en3, QN => n_1404);
   cw2_reg_6_inst : DLH_X1 port map( G => N174, D => n91, Q => cw2_6_port);
   cw3_reg_6_inst : SDFF_X1 port map( D => n14, SI => n85, SE => cw2_6_port, CK
                           => Clk, Q => Mux1Sel, QN => n_1405);
   cw2_reg_5_inst : DLH_X1 port map( G => N174, D => n88, Q => cw2_5_port);
   cw2_reg_4_inst : DLH_X1 port map( G => N174, D => n85, Q => cw2_4_port);
   cw3_reg_4_inst : SDFF_X1 port map( D => n12, SI => n85, SE => cw2_4_port, CK
                           => Clk, Q => n_1406, QN => n362);
   cw2_reg_3_inst : DLH_X1 port map( G => N174, D => n94, Q => cw2_3_port);
   cw3_reg_3_inst : SDFF_X1 port map( D => n10, SI => n85, SE => cw2_3_port, CK
                           => Clk, Q => n_1407, QN => n361);
   cw2_reg_2_inst : DLH_X1 port map( G => N174, D => N176, Q => cw2_2_port);
   cw3_reg_2_inst : SDFF_X1 port map( D => n8, SI => n85, SE => cw2_2_port, CK 
                           => Clk, Q => n_1408, QN => n360);
   cw2_reg_1_inst : DLH_X1 port map( G => N174, D => N176, Q => cw2_1_port);
   cw3_reg_1_inst : SDFF_X1 port map( D => n6, SI => n85, SE => cw2_1_port, CK 
                           => Clk, Q => n_1409, QN => n359);
   cw2_reg_0_inst : DLH_X1 port map( G => N174, D => N175, Q => cw2_0_port);
   cw3_reg_0_inst : SDFF_X1 port map( D => n3, SI => n85, SE => cw2_0_port, CK 
                           => Clk, Q => n_1410, QN => n358);
   n3 <= '0';
   n6 <= '0';
   n8 <= '0';
   n10 <= '0';
   n12 <= '0';
   n13 <= '0';
   n14 <= '0';
   n15 <= '0';
   cw5_reg_0_inst : DFF_X1 port map( D => n282, CK => Clk, Q => WR, QN => 
                           n_1411);
   cw4_reg_4_inst : DFF_X1 port map( D => n281, CK => Clk, Q => en4, QN => 
                           n_1412);
   cw4_reg_3_inst : DFF_X1 port map( D => n280, CK => Clk, Q => MemoryEnable, 
                           QN => n_1413);
   cw4_reg_2_inst : DFF_X1 port map( D => n279, CK => Clk, Q => ReadNotWrite, 
                           QN => n_1414);
   cw4_reg_1_inst : DFF_X1 port map( D => n278, CK => Clk, Q => n_1415, QN => 
                           n275);
   cw4_reg_0_inst : DFF_X1 port map( D => n277, CK => Clk, Q => n_1416, QN => 
                           n276);
   U296 : OAI33_X1 port map( A1 => n111, A2 => n317, A3 => n318, B1 => n319, B2
                           => n320, B3 => n321, ZN => n316);
   U297 : NAND3_X1 port map( A1 => n86, A2 => n320, A3 => n107, ZN => n331);
   U298 : NAND3_X1 port map( A1 => n352, A2 => n349, A3 => n353, ZN => N174);
   U299 : NAND3_X1 port map( A1 => IR_IN(28), A2 => n354, A3 => IR_IN(30), ZN 
                           => n327);
   U300 : NAND3_X1 port map( A1 => n365, A2 => n96, A3 => n340, ZN => n332);
   U301 : NAND3_X1 port map( A1 => n366, A2 => n98, A3 => n326, ZN => n365);
   U302 : NAND3_X1 port map( A1 => n340, A2 => n367, A3 => IR_IN(30), ZN => 
                           n330);
   U303 : NAND3_X1 port map( A1 => IR_IN(26), A2 => n355, A3 => IR_IN(31), ZN 
                           => n342);
   cw3_reg_5_inst : SDFF_X1 port map( D => n13, SI => n85, SE => cw2_5_port, CK
                           => Clk, Q => Mux2Sel, QN => n_1417);
   cw2_reg_14_inst : DLH_X1 port map( G => N174, D => N185, Q => SignSelect);
   cw5_reg_1_inst : DFF_X1 port map( D => n283, CK => Clk, Q => selwb, QN => 
                           n_1418);
   aluOpcode3_reg_0_inst : DFF_X1 port map( D => n103, CK => Clk, Q => 
                           ALUCODE_0_port, QN => n193);
   U210 : INV_X1 port map( A => n318, ZN => n88);
   U211 : INV_X1 port map( A => n321, ZN => n106);
   U212 : INV_X1 port map( A => n319, ZN => n86);
   U213 : NAND2_X1 port map( A1 => n329, A2 => n318, ZN => N183);
   U214 : OR2_X1 port map( A1 => n88, A2 => N185, ZN => N184);
   U215 : INV_X1 port map( A => n313, ZN => n90);
   U216 : INV_X1 port map( A => n329, ZN => n94);
   U217 : NAND4_X1 port map( A1 => n340, A2 => n341, A3 => n99, A4 => n96, ZN 
                           => n343);
   U218 : NAND4_X1 port map( A1 => n110, A2 => n109, A3 => n108, A4 => n339, ZN
                           => n324);
   U219 : NAND2_X1 port map( A1 => n348, A2 => n85, ZN => n318);
   U220 : NAND2_X1 port map( A1 => n338, A2 => n110, ZN => n321);
   U221 : AND3_X1 port map( A1 => n351, A2 => n99, A3 => n341, ZN => n348);
   U222 : AND2_X1 port map( A1 => n354, A2 => n96, ZN => n351);
   U223 : AND2_X1 port map( A1 => n354, A2 => n355, ZN => n346);
   U224 : INV_X1 port map( A => n366, ZN => n100);
   U225 : INV_X1 port map( A => n340, ZN => n93);
   U226 : INV_X1 port map( A => n327, ZN => n92);
   U227 : NAND2_X1 port map( A1 => n88, A2 => n112, ZN => n319);
   U228 : INV_X1 port map( A => n356, ZN => n98);
   U229 : INV_X1 port map( A => n328, ZN => n89);
   U230 : NAND2_X1 port map( A1 => n111, A2 => n113, ZN => n320);
   U231 : AOI21_X1 port map( B1 => n100, B2 => n351, A => n95, ZN => n352);
   U232 : NOR4_X1 port map( A1 => Rst, A2 => n348, A3 => n350, A4 => n346, ZN 
                           => n353);
   U233 : AOI21_X1 port map( B1 => n85, B2 => n350, A => n364, ZN => n313);
   U234 : NAND2_X1 port map( A1 => n95, A2 => n85, ZN => n329);
   U235 : OAI211_X1 port map( C1 => Rst, C2 => n349, A => n329, B => n313, ZN 
                           => N185);
   U236 : INV_X1 port map( A => n342, ZN => n95);
   U237 : OAI211_X1 port map( C1 => Rst, C2 => n349, A => n318, B => n312, ZN 
                           => N175);
   U238 : AND2_X1 port map( A1 => n356, A2 => n351, ZN => n350);
   U239 : AND3_X1 port map( A1 => n351, A2 => n85, A3 => n100, ZN => n364);
   U240 : AND2_X1 port map( A1 => n346, A2 => n85, ZN => N182);
   U241 : INV_X1 port map( A => n312, ZN => n91);
   U242 : NOR4_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), A3 => IR_IN(7), A4 
                           => IR_IN(6), ZN => n339);
   U243 : INV_X1 port map( A => n314, ZN => n87);
   U244 : AOI221_X1 port map( B1 => n315, B2 => n85, C1 => Rst, C2 => 
                           ALUCODE_1_port, A => n316, ZN => n314);
   U245 : OAI221_X1 port map( B1 => n98, B2 => n93, C1 => n326, C2 => n327, A 
                           => n89, ZN => n315);
   U246 : NOR2_X1 port map( A1 => n97, A2 => IR_IN(31), ZN => n340);
   U247 : NOR2_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), ZN => n341);
   U248 : NOR3_X1 port map( A1 => n101, A2 => IR_IN(27), A3 => n99, ZN => n356)
                           ;
   U249 : NOR2_X1 port map( A1 => n112, A2 => IR_IN(0), ZN => n323);
   U250 : OAI221_X1 port map( B1 => Rst, B2 => n335, C1 => n193, C2 => n85, A 
                           => n336, ZN => n103);
   U251 : OAI211_X1 port map( C1 => n337, C2 => n106, A => n113, B => n86, ZN 
                           => n336);
   U252 : AOI221_X1 port map( B1 => n340, B2 => n100, C1 => n92, C2 => n341, A 
                           => n328, ZN => n335);
   U253 : AOI21_X1 port map( B1 => n324, B2 => n325, A => n111, ZN => n337);
   U254 : NAND2_X1 port map( A1 => IR_IN(27), A2 => n101, ZN => n326);
   U255 : NAND4_X1 port map( A1 => n342, A2 => n343, A3 => n344, A4 => n345, ZN
                           => n328);
   U256 : AOI21_X1 port map( B1 => IR_IN(26), B2 => n346, A => n347, ZN => n345
                           );
   U257 : NAND4_X1 port map( A1 => IR_IN(2), A2 => n323, A3 => n106, A4 => n348
                           , ZN => n344);
   U258 : NOR4_X1 port map( A1 => IR_IN(30), A2 => n99, A3 => n93, A4 => n326, 
                           ZN => n347);
   U259 : NOR2_X1 port map( A1 => IR_IN(29), A2 => IR_IN(31), ZN => n354);
   U260 : AOI22_X1 port map( A1 => n322, A2 => IR_IN(0), B1 => n323, B2 => n102
                           , ZN => n317);
   U261 : INV_X1 port map( A => n324, ZN => n102);
   U262 : AOI21_X1 port map( B1 => n321, B2 => n325, A => IR_IN(1), ZN => n322)
                           ;
   U263 : INV_X1 port map( A => IR_IN(28), ZN => n99);
   U264 : NAND2_X1 port map( A1 => IR_IN(3), A2 => n338, ZN => n325);
   U265 : NAND2_X1 port map( A1 => n341, A2 => IR_IN(28), ZN => n366);
   U266 : OAI21_X1 port map( B1 => IR_IN(27), B2 => n101, A => n366, ZN => n367
                           );
   U267 : INV_X1 port map( A => IR_IN(26), ZN => n101);
   U268 : OAI221_X1 port map( B1 => Rst, B2 => n330, C1 => n195, C2 => n85, A 
                           => n331, ZN => n105);
   U269 : INV_X1 port map( A => n325, ZN => n107);
   U270 : INV_X1 port map( A => IR_IN(1), ZN => n112);
   U271 : INV_X1 port map( A => IR_IN(30), ZN => n96);
   U272 : INV_X1 port map( A => IR_IN(2), ZN => n111);
   U273 : INV_X1 port map( A => IR_IN(0), ZN => n113);
   U274 : AND4_X1 port map( A1 => n108, A2 => n109, A3 => IR_IN(5), A4 => n339,
                           ZN => n338);
   U275 : INV_X1 port map( A => IR_IN(3), ZN => n110);
   U276 : INV_X1 port map( A => IR_IN(29), ZN => n97);
   U277 : INV_X1 port map( A => IR_IN(4), ZN => n109);
   U278 : INV_X1 port map( A => IR_IN(10), ZN => n108);
   U279 : AND3_X1 port map( A1 => n99, A2 => n96, A3 => IR_IN(27), ZN => n355);
   U280 : OAI221_X1 port map( B1 => Rst, B2 => n332, C1 => n194, C2 => n85, A 
                           => n333, ZN => n104);
   U281 : OR3_X1 port map( A1 => n318, A2 => n334, A3 => n321, ZN => n333);
   U282 : AOI21_X1 port map( B1 => n112, B2 => IR_IN(2), A => n323, ZN => n334)
                           ;
   U283 : NOR2_X1 port map( A1 => Rst, A2 => n358, ZN => n277);
   U284 : NOR2_X1 port map( A1 => Rst, A2 => n359, ZN => n278);
   U285 : NOR2_X1 port map( A1 => Rst, A2 => n360, ZN => n279);
   U286 : NOR2_X1 port map( A1 => Rst, A2 => n361, ZN => n280);
   U287 : NOR2_X1 port map( A1 => Rst, A2 => n362, ZN => n281);
   U288 : NOR2_X1 port map( A1 => Rst, A2 => n276, ZN => n282);
   U289 : NOR2_X1 port map( A1 => Rst, A2 => n275, ZN => n283);
   U290 : INV_X1 port map( A => Rst, ZN => n85);
   U291 : NAND2_X1 port map( A1 => IR_IN(26), A2 => N182, ZN => n312);
   U292 : NOR2_X1 port map( A1 => IR_IN(29), A2 => n329, ZN => N176);
   U293 : AND4_X1 port map( A1 => n330, A2 => n343, A3 => n332, A4 => n357, ZN 
                           => n349);
   U294 : AOI21_X1 port map( B1 => n95, B2 => n97, A => n363, ZN => n357);
   U295 : AOI21_X1 port map( B1 => IR_IN(27), B2 => n326, A => n327, ZN => n363
                           );

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_M32_C4_N5.all;

entity DLX_M32_C4_N5 is

   port( Clk, Rst : in std_logic;  IRAM_Addr : out std_logic_vector (31 downto 
         0);  IRAM_Dout : in std_logic_vector (31 downto 0);  DRAM_MemoryEnable
         , DRAM_ReadNotWrite : out std_logic;  DRAM_Addr : out std_logic_vector
         (4 downto 0);  DRAM_in : out std_logic_vector (31 downto 0);  DRAM_out
         : in std_logic_vector (31 downto 0));

end DLX_M32_C4_N5;

architecture SYN_dlx_rtl of DLX_M32_C4_N5 is

   component dataPath_M32_C4_N5
      port( clock, reset : in std_logic;  Instruction : in std_logic_vector (31
            downto 0);  en1, en2, SignSelect, RD1, RD2, WR, JMP, BRANCHenable, 
            en3, BranchCondSel, Mux1Sel, Mux2Sel : in std_logic;  ALUCODE : in 
            std_logic_vector (3 downto 0);  RegDestination, en4 : in std_logic;
            DRAMout : in std_logic_vector (31 downto 0);  selwb : in std_logic;
            PCtoIM, ALUtoMEMORY, OUT2RFtoMEMORY, InstructionToCU : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  en1, en2, SignSelect, RD1, RD2, JMP, BranchCondSel, BRANCHenable
            , RegDestination, en3, Mux1Sel, Mux2Sel : out std_logic;  ALUCODE :
            out std_logic_vector (3 downto 0);  en4, MemoryEnable, ReadNotWrite
            , selwb, WR : out std_logic);
   end component;
   
   signal InstructionToCU_31_port, InstructionToCU_30_port, 
      InstructionToCU_29_port, InstructionToCU_28_port, InstructionToCU_27_port
      , InstructionToCU_26_port, InstructionToCU_25_port, 
      InstructionToCU_24_port, InstructionToCU_23_port, InstructionToCU_22_port
      , InstructionToCU_21_port, InstructionToCU_20_port, 
      InstructionToCU_19_port, InstructionToCU_18_port, InstructionToCU_17_port
      , InstructionToCU_16_port, InstructionToCU_15_port, 
      InstructionToCU_14_port, InstructionToCU_13_port, InstructionToCU_12_port
      , InstructionToCU_11_port, InstructionToCU_10_port, 
      InstructionToCU_9_port, InstructionToCU_8_port, InstructionToCU_7_port, 
      InstructionToCU_6_port, InstructionToCU_5_port, InstructionToCU_4_port, 
      InstructionToCU_3_port, InstructionToCU_2_port, InstructionToCU_1_port, 
      InstructionToCU_0_port, en1, en2, SignSelect, RD1, RD2, JMP, 
      BranchCondSel, BRANCHenable, RegDestination, en3, Mux1Sel, Mux2Sel, 
      ALUCODE_3_port, ALUCODE_2_port, ALUCODE_1_port, ALUCODE_0_port, en4, 
      selwb, WR, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426
      , n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435,
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446 : std_logic;

begin
   
   en1 <= '1';
   CU_I : Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17 port 
                           map( Clk => Clk, Rst => Rst, IR_IN(31) => 
                           InstructionToCU_31_port, IR_IN(30) => 
                           InstructionToCU_30_port, IR_IN(29) => 
                           InstructionToCU_29_port, IR_IN(28) => 
                           InstructionToCU_28_port, IR_IN(27) => 
                           InstructionToCU_27_port, IR_IN(26) => 
                           InstructionToCU_26_port, IR_IN(25) => 
                           InstructionToCU_25_port, IR_IN(24) => 
                           InstructionToCU_24_port, IR_IN(23) => 
                           InstructionToCU_23_port, IR_IN(22) => 
                           InstructionToCU_22_port, IR_IN(21) => 
                           InstructionToCU_21_port, IR_IN(20) => 
                           InstructionToCU_20_port, IR_IN(19) => 
                           InstructionToCU_19_port, IR_IN(18) => 
                           InstructionToCU_18_port, IR_IN(17) => 
                           InstructionToCU_17_port, IR_IN(16) => 
                           InstructionToCU_16_port, IR_IN(15) => 
                           InstructionToCU_15_port, IR_IN(14) => 
                           InstructionToCU_14_port, IR_IN(13) => 
                           InstructionToCU_13_port, IR_IN(12) => 
                           InstructionToCU_12_port, IR_IN(11) => 
                           InstructionToCU_11_port, IR_IN(10) => 
                           InstructionToCU_10_port, IR_IN(9) => 
                           InstructionToCU_9_port, IR_IN(8) => 
                           InstructionToCU_8_port, IR_IN(7) => 
                           InstructionToCU_7_port, IR_IN(6) => 
                           InstructionToCU_6_port, IR_IN(5) => 
                           InstructionToCU_5_port, IR_IN(4) => 
                           InstructionToCU_4_port, IR_IN(3) => 
                           InstructionToCU_3_port, IR_IN(2) => 
                           InstructionToCU_2_port, IR_IN(1) => 
                           InstructionToCU_1_port, IR_IN(0) => 
                           InstructionToCU_0_port, en1 => n_1419, en2 => en2, 
                           SignSelect => SignSelect, RD1 => RD1, RD2 => RD2, 
                           JMP => JMP, BranchCondSel => BranchCondSel, 
                           BRANCHenable => BRANCHenable, RegDestination => 
                           RegDestination, en3 => en3, Mux1Sel => Mux1Sel, 
                           Mux2Sel => Mux2Sel, ALUCODE(3) => ALUCODE_3_port, 
                           ALUCODE(2) => ALUCODE_2_port, ALUCODE(1) => 
                           ALUCODE_1_port, ALUCODE(0) => ALUCODE_0_port, en4 =>
                           en4, MemoryEnable => DRAM_MemoryEnable, ReadNotWrite
                           => DRAM_ReadNotWrite, selwb => selwb, WR => WR);
   DP : dataPath_M32_C4_N5 port map( clock => Clk, reset => Rst, 
                           Instruction(31) => IRAM_Dout(31), Instruction(30) =>
                           IRAM_Dout(30), Instruction(29) => IRAM_Dout(29), 
                           Instruction(28) => IRAM_Dout(28), Instruction(27) =>
                           IRAM_Dout(27), Instruction(26) => IRAM_Dout(26), 
                           Instruction(25) => IRAM_Dout(25), Instruction(24) =>
                           IRAM_Dout(24), Instruction(23) => IRAM_Dout(23), 
                           Instruction(22) => IRAM_Dout(22), Instruction(21) =>
                           IRAM_Dout(21), Instruction(20) => IRAM_Dout(20), 
                           Instruction(19) => IRAM_Dout(19), Instruction(18) =>
                           IRAM_Dout(18), Instruction(17) => IRAM_Dout(17), 
                           Instruction(16) => IRAM_Dout(16), Instruction(15) =>
                           IRAM_Dout(15), Instruction(14) => IRAM_Dout(14), 
                           Instruction(13) => IRAM_Dout(13), Instruction(12) =>
                           IRAM_Dout(12), Instruction(11) => IRAM_Dout(11), 
                           Instruction(10) => IRAM_Dout(10), Instruction(9) => 
                           IRAM_Dout(9), Instruction(8) => IRAM_Dout(8), 
                           Instruction(7) => IRAM_Dout(7), Instruction(6) => 
                           IRAM_Dout(6), Instruction(5) => IRAM_Dout(5), 
                           Instruction(4) => IRAM_Dout(4), Instruction(3) => 
                           IRAM_Dout(3), Instruction(2) => IRAM_Dout(2), 
                           Instruction(1) => IRAM_Dout(1), Instruction(0) => 
                           IRAM_Dout(0), en1 => en1, en2 => en2, SignSelect => 
                           SignSelect, RD1 => RD1, RD2 => RD2, WR => WR, JMP =>
                           JMP, BRANCHenable => BRANCHenable, en3 => en3, 
                           BranchCondSel => BranchCondSel, Mux1Sel => Mux1Sel, 
                           Mux2Sel => Mux2Sel, ALUCODE(3) => ALUCODE_3_port, 
                           ALUCODE(2) => ALUCODE_2_port, ALUCODE(1) => 
                           ALUCODE_1_port, ALUCODE(0) => ALUCODE_0_port, 
                           RegDestination => RegDestination, en4 => en4, 
                           DRAMout(31) => DRAM_out(31), DRAMout(30) => 
                           DRAM_out(30), DRAMout(29) => DRAM_out(29), 
                           DRAMout(28) => DRAM_out(28), DRAMout(27) => 
                           DRAM_out(27), DRAMout(26) => DRAM_out(26), 
                           DRAMout(25) => DRAM_out(25), DRAMout(24) => 
                           DRAM_out(24), DRAMout(23) => DRAM_out(23), 
                           DRAMout(22) => DRAM_out(22), DRAMout(21) => 
                           DRAM_out(21), DRAMout(20) => DRAM_out(20), 
                           DRAMout(19) => DRAM_out(19), DRAMout(18) => 
                           DRAM_out(18), DRAMout(17) => DRAM_out(17), 
                           DRAMout(16) => DRAM_out(16), DRAMout(15) => 
                           DRAM_out(15), DRAMout(14) => DRAM_out(14), 
                           DRAMout(13) => DRAM_out(13), DRAMout(12) => 
                           DRAM_out(12), DRAMout(11) => DRAM_out(11), 
                           DRAMout(10) => DRAM_out(10), DRAMout(9) => 
                           DRAM_out(9), DRAMout(8) => DRAM_out(8), DRAMout(7) 
                           => DRAM_out(7), DRAMout(6) => DRAM_out(6), 
                           DRAMout(5) => DRAM_out(5), DRAMout(4) => DRAM_out(4)
                           , DRAMout(3) => DRAM_out(3), DRAMout(2) => 
                           DRAM_out(2), DRAMout(1) => DRAM_out(1), DRAMout(0) 
                           => DRAM_out(0), selwb => selwb, PCtoIM(31) => 
                           IRAM_Addr(31), PCtoIM(30) => IRAM_Addr(30), 
                           PCtoIM(29) => IRAM_Addr(29), PCtoIM(28) => 
                           IRAM_Addr(28), PCtoIM(27) => IRAM_Addr(27), 
                           PCtoIM(26) => IRAM_Addr(26), PCtoIM(25) => 
                           IRAM_Addr(25), PCtoIM(24) => IRAM_Addr(24), 
                           PCtoIM(23) => IRAM_Addr(23), PCtoIM(22) => 
                           IRAM_Addr(22), PCtoIM(21) => IRAM_Addr(21), 
                           PCtoIM(20) => IRAM_Addr(20), PCtoIM(19) => 
                           IRAM_Addr(19), PCtoIM(18) => IRAM_Addr(18), 
                           PCtoIM(17) => IRAM_Addr(17), PCtoIM(16) => 
                           IRAM_Addr(16), PCtoIM(15) => IRAM_Addr(15), 
                           PCtoIM(14) => IRAM_Addr(14), PCtoIM(13) => 
                           IRAM_Addr(13), PCtoIM(12) => IRAM_Addr(12), 
                           PCtoIM(11) => IRAM_Addr(11), PCtoIM(10) => 
                           IRAM_Addr(10), PCtoIM(9) => IRAM_Addr(9), PCtoIM(8) 
                           => IRAM_Addr(8), PCtoIM(7) => IRAM_Addr(7), 
                           PCtoIM(6) => IRAM_Addr(6), PCtoIM(5) => IRAM_Addr(5)
                           , PCtoIM(4) => IRAM_Addr(4), PCtoIM(3) => 
                           IRAM_Addr(3), PCtoIM(2) => IRAM_Addr(2), PCtoIM(1) 
                           => IRAM_Addr(1), PCtoIM(0) => IRAM_Addr(0), 
                           ALUtoMEMORY(31) => n_1420, ALUtoMEMORY(30) => n_1421
                           , ALUtoMEMORY(29) => n_1422, ALUtoMEMORY(28) => 
                           n_1423, ALUtoMEMORY(27) => n_1424, ALUtoMEMORY(26) 
                           => n_1425, ALUtoMEMORY(25) => n_1426, 
                           ALUtoMEMORY(24) => n_1427, ALUtoMEMORY(23) => n_1428
                           , ALUtoMEMORY(22) => n_1429, ALUtoMEMORY(21) => 
                           n_1430, ALUtoMEMORY(20) => n_1431, ALUtoMEMORY(19) 
                           => n_1432, ALUtoMEMORY(18) => n_1433, 
                           ALUtoMEMORY(17) => n_1434, ALUtoMEMORY(16) => n_1435
                           , ALUtoMEMORY(15) => n_1436, ALUtoMEMORY(14) => 
                           n_1437, ALUtoMEMORY(13) => n_1438, ALUtoMEMORY(12) 
                           => n_1439, ALUtoMEMORY(11) => n_1440, 
                           ALUtoMEMORY(10) => n_1441, ALUtoMEMORY(9) => n_1442,
                           ALUtoMEMORY(8) => n_1443, ALUtoMEMORY(7) => n_1444, 
                           ALUtoMEMORY(6) => n_1445, ALUtoMEMORY(5) => n_1446, 
                           ALUtoMEMORY(4) => DRAM_Addr(4), ALUtoMEMORY(3) => 
                           DRAM_Addr(3), ALUtoMEMORY(2) => DRAM_Addr(2), 
                           ALUtoMEMORY(1) => DRAM_Addr(1), ALUtoMEMORY(0) => 
                           DRAM_Addr(0), OUT2RFtoMEMORY(31) => DRAM_in(31), 
                           OUT2RFtoMEMORY(30) => DRAM_in(30), 
                           OUT2RFtoMEMORY(29) => DRAM_in(29), 
                           OUT2RFtoMEMORY(28) => DRAM_in(28), 
                           OUT2RFtoMEMORY(27) => DRAM_in(27), 
                           OUT2RFtoMEMORY(26) => DRAM_in(26), 
                           OUT2RFtoMEMORY(25) => DRAM_in(25), 
                           OUT2RFtoMEMORY(24) => DRAM_in(24), 
                           OUT2RFtoMEMORY(23) => DRAM_in(23), 
                           OUT2RFtoMEMORY(22) => DRAM_in(22), 
                           OUT2RFtoMEMORY(21) => DRAM_in(21), 
                           OUT2RFtoMEMORY(20) => DRAM_in(20), 
                           OUT2RFtoMEMORY(19) => DRAM_in(19), 
                           OUT2RFtoMEMORY(18) => DRAM_in(18), 
                           OUT2RFtoMEMORY(17) => DRAM_in(17), 
                           OUT2RFtoMEMORY(16) => DRAM_in(16), 
                           OUT2RFtoMEMORY(15) => DRAM_in(15), 
                           OUT2RFtoMEMORY(14) => DRAM_in(14), 
                           OUT2RFtoMEMORY(13) => DRAM_in(13), 
                           OUT2RFtoMEMORY(12) => DRAM_in(12), 
                           OUT2RFtoMEMORY(11) => DRAM_in(11), 
                           OUT2RFtoMEMORY(10) => DRAM_in(10), OUT2RFtoMEMORY(9)
                           => DRAM_in(9), OUT2RFtoMEMORY(8) => DRAM_in(8), 
                           OUT2RFtoMEMORY(7) => DRAM_in(7), OUT2RFtoMEMORY(6) 
                           => DRAM_in(6), OUT2RFtoMEMORY(5) => DRAM_in(5), 
                           OUT2RFtoMEMORY(4) => DRAM_in(4), OUT2RFtoMEMORY(3) 
                           => DRAM_in(3), OUT2RFtoMEMORY(2) => DRAM_in(2), 
                           OUT2RFtoMEMORY(1) => DRAM_in(1), OUT2RFtoMEMORY(0) 
                           => DRAM_in(0), InstructionToCU(31) => 
                           InstructionToCU_31_port, InstructionToCU(30) => 
                           InstructionToCU_30_port, InstructionToCU(29) => 
                           InstructionToCU_29_port, InstructionToCU(28) => 
                           InstructionToCU_28_port, InstructionToCU(27) => 
                           InstructionToCU_27_port, InstructionToCU(26) => 
                           InstructionToCU_26_port, InstructionToCU(25) => 
                           InstructionToCU_25_port, InstructionToCU(24) => 
                           InstructionToCU_24_port, InstructionToCU(23) => 
                           InstructionToCU_23_port, InstructionToCU(22) => 
                           InstructionToCU_22_port, InstructionToCU(21) => 
                           InstructionToCU_21_port, InstructionToCU(20) => 
                           InstructionToCU_20_port, InstructionToCU(19) => 
                           InstructionToCU_19_port, InstructionToCU(18) => 
                           InstructionToCU_18_port, InstructionToCU(17) => 
                           InstructionToCU_17_port, InstructionToCU(16) => 
                           InstructionToCU_16_port, InstructionToCU(15) => 
                           InstructionToCU_15_port, InstructionToCU(14) => 
                           InstructionToCU_14_port, InstructionToCU(13) => 
                           InstructionToCU_13_port, InstructionToCU(12) => 
                           InstructionToCU_12_port, InstructionToCU(11) => 
                           InstructionToCU_11_port, InstructionToCU(10) => 
                           InstructionToCU_10_port, InstructionToCU(9) => 
                           InstructionToCU_9_port, InstructionToCU(8) => 
                           InstructionToCU_8_port, InstructionToCU(7) => 
                           InstructionToCU_7_port, InstructionToCU(6) => 
                           InstructionToCU_6_port, InstructionToCU(5) => 
                           InstructionToCU_5_port, InstructionToCU(4) => 
                           InstructionToCU_4_port, InstructionToCU(3) => 
                           InstructionToCU_3_port, InstructionToCU(2) => 
                           InstructionToCU_2_port, InstructionToCU(1) => 
                           InstructionToCU_1_port, InstructionToCU(0) => 
                           InstructionToCU_0_port);

end SYN_dlx_rtl;
