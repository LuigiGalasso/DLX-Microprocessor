
module Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17 ( Clk, Rst, 
        IR_IN, en1, en2, SignSelect, RD1, RD2, JMP, BranchCondSel, 
        BRANCHenable, RegDestination, en3, Mux1Sel, Mux2Sel, ALUCODE, en4, 
        MemoryEnable, ReadNotWrite, selwb, WR );
  input [31:0] IR_IN;
  output [3:0] ALUCODE;
  input Clk, Rst;
  output en1, en2, SignSelect, RD1, RD2, JMP, BranchCondSel, BRANCHenable,
         RegDestination, en3, Mux1Sel, Mux2Sel, en4, MemoryEnable,
         ReadNotWrite, selwb, WR;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26, N174,
         N175, N176, N182, N183, N184, N185, n103, n104, n105, n193, n194,
         n195, n275, n276, n277, n278, n279, n280, n281, n282, n283, n358,
         n359, n360, n361, n362, n364, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n363, n365, n366, n367, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n106, n107, n108, n109, n110, n111, n112;
  wire   [7:0] cw2;
  assign en1 = 1'b1;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];

  DFF_X1 \aluOpcode3_reg[3]  ( .D(n105), .CK(Clk), .Q(ALUCODE[3]), .QN(n195)
         );
  DFF_X1 \aluOpcode3_reg[2]  ( .D(n104), .CK(Clk), .Q(ALUCODE[2]), .QN(n194)
         );
  DFF_X1 \aluOpcode3_reg[1]  ( .D(n85), .CK(Clk), .Q(ALUCODE[1]) );
  DLH_X1 \cw2_reg[15]  ( .G(N174), .D(n84), .Q(en2) );
  DLH_X1 \cw2_reg[14]  ( .G(N174), .D(N185), .Q(SignSelect) );
  DLH_X1 \cw2_reg[13]  ( .G(N174), .D(N184), .Q(RD1) );
  DLH_X1 \cw2_reg[12]  ( .G(N174), .D(N183), .Q(RD2) );
  DLH_X1 \cw2_reg[11]  ( .G(N174), .D(N182), .Q(JMP) );
  DLH_X1 \cw2_reg[10]  ( .G(N174), .D(n364), .Q(BranchCondSel) );
  DLH_X1 \cw2_reg[9]  ( .G(N174), .D(n90), .Q(BRANCHenable) );
  DLH_X1 \cw2_reg[8]  ( .G(N174), .D(n88), .Q(RegDestination) );
  DLH_X1 \cw2_reg[7]  ( .G(N174), .D(n84), .Q(cw2[7]) );
  SDFF_X1 \cw3_reg[7]  ( .D(1'b0), .SI(n84), .SE(cw2[7]), .CK(Clk), .Q(en3) );
  DLH_X1 \cw2_reg[6]  ( .G(N174), .D(n91), .Q(cw2[6]) );
  SDFF_X1 \cw3_reg[6]  ( .D(1'b0), .SI(n84), .SE(cw2[6]), .CK(Clk), .Q(Mux1Sel) );
  DLH_X1 \cw2_reg[5]  ( .G(N174), .D(n88), .Q(cw2[5]) );
  DLH_X1 \cw2_reg[4]  ( .G(N174), .D(n84), .Q(cw2[4]) );
  SDFF_X1 \cw3_reg[4]  ( .D(1'b0), .SI(n84), .SE(cw2[4]), .CK(Clk), .QN(n362)
         );
  DLH_X1 \cw2_reg[3]  ( .G(N174), .D(n92), .Q(cw2[3]) );
  SDFF_X1 \cw3_reg[3]  ( .D(1'b0), .SI(n84), .SE(cw2[3]), .CK(Clk), .QN(n361)
         );
  DLH_X1 \cw2_reg[2]  ( .G(N174), .D(N176), .Q(cw2[2]) );
  SDFF_X1 \cw3_reg[2]  ( .D(1'b0), .SI(n84), .SE(cw2[2]), .CK(Clk), .QN(n360)
         );
  DLH_X1 \cw2_reg[1]  ( .G(N174), .D(N176), .Q(cw2[1]) );
  SDFF_X1 \cw3_reg[1]  ( .D(1'b0), .SI(n84), .SE(cw2[1]), .CK(Clk), .QN(n359)
         );
  DLH_X1 \cw2_reg[0]  ( .G(N174), .D(N175), .Q(cw2[0]) );
  SDFF_X1 \cw3_reg[0]  ( .D(1'b0), .SI(n84), .SE(cw2[0]), .CK(Clk), .QN(n358)
         );
  DFF_X1 \cw5_reg[0]  ( .D(n282), .CK(Clk), .Q(WR) );
  DFF_X1 \cw4_reg[4]  ( .D(n281), .CK(Clk), .Q(en4) );
  DFF_X1 \cw4_reg[3]  ( .D(n280), .CK(Clk), .Q(MemoryEnable) );
  DFF_X1 \cw4_reg[2]  ( .D(n279), .CK(Clk), .Q(ReadNotWrite) );
  DFF_X1 \cw4_reg[1]  ( .D(n278), .CK(Clk), .QN(n275) );
  DFF_X1 \cw4_reg[0]  ( .D(n277), .CK(Clk), .QN(n276) );
  OAI33_X1 U296 ( .A1(n110), .A2(n318), .A3(n319), .B1(n320), .B2(n321), .B3(
        n322), .ZN(n317) );
  NAND3_X1 U297 ( .A1(n87), .A2(n321), .A3(n100), .ZN(n331) );
  NAND3_X1 U298 ( .A1(n352), .A2(n349), .A3(n353), .ZN(N174) );
  NAND3_X1 U299 ( .A1(n355), .A2(IR_IN_28), .A3(IR_IN_30), .ZN(n328) );
  NAND3_X1 U300 ( .A1(n365), .A2(n98), .A3(n340), .ZN(n332) );
  NAND3_X1 U301 ( .A1(n89), .A2(n327), .A3(n366), .ZN(n365) );
  NAND3_X1 U302 ( .A1(n340), .A2(n367), .A3(IR_IN_30), .ZN(n330) );
  NAND3_X1 U303 ( .A1(n354), .A2(IR_IN_26), .A3(IR_IN_31), .ZN(n342) );
  SDFF_X1 \cw3_reg[5]  ( .D(1'b0), .SI(n84), .SE(cw2[5]), .CK(Clk), .Q(Mux2Sel) );
  DFF_X1 \aluOpcode3_reg[0]  ( .D(n103), .CK(Clk), .Q(ALUCODE[0]), .QN(n193)
         );
  DFF_X1 \cw5_reg[1]  ( .D(n283), .CK(Clk), .Q(selwb) );
  INV_X1 U210 ( .A(n319), .ZN(n88) );
  INV_X1 U211 ( .A(n322), .ZN(n99) );
  INV_X1 U212 ( .A(n320), .ZN(n87) );
  NAND2_X1 U213 ( .A1(n314), .A2(n319), .ZN(N183) );
  OR2_X1 U214 ( .A1(n88), .A2(N185), .ZN(N184) );
  INV_X1 U215 ( .A(n312), .ZN(n90) );
  INV_X1 U216 ( .A(n314), .ZN(n92) );
  NAND4_X1 U217 ( .A1(n340), .A2(n341), .A3(n94), .A4(n98), .ZN(n343) );
  NAND4_X1 U218 ( .A1(n107), .A2(n106), .A3(n102), .A4(n339), .ZN(n325) );
  NAND2_X1 U219 ( .A1(n348), .A2(n84), .ZN(n319) );
  NAND2_X1 U220 ( .A1(n338), .A2(n107), .ZN(n322) );
  AND3_X1 U221 ( .A1(n351), .A2(n94), .A3(n341), .ZN(n348) );
  AND2_X1 U222 ( .A1(n355), .A2(n98), .ZN(n351) );
  AND2_X1 U223 ( .A1(n354), .A2(n355), .ZN(n346) );
  INV_X1 U224 ( .A(n366), .ZN(n95) );
  INV_X1 U225 ( .A(n340), .ZN(n109) );
  INV_X1 U226 ( .A(n328), .ZN(n96) );
  NAND2_X1 U227 ( .A1(n88), .A2(n108), .ZN(n320) );
  INV_X1 U228 ( .A(n356), .ZN(n89) );
  INV_X1 U229 ( .A(n329), .ZN(n86) );
  NAND2_X1 U230 ( .A1(n110), .A2(n111), .ZN(n321) );
  AOI21_X1 U231 ( .B1(n95), .B2(n351), .A(n93), .ZN(n352) );
  NOR4_X1 U232 ( .A1(Rst), .A2(n350), .A3(n348), .A4(n346), .ZN(n353) );
  AOI21_X1 U233 ( .B1(n84), .B2(n350), .A(n364), .ZN(n312) );
  NAND2_X1 U234 ( .A1(n93), .A2(n84), .ZN(n314) );
  OAI211_X1 U235 ( .C1(Rst), .C2(n349), .A(n314), .B(n312), .ZN(N185) );
  INV_X1 U236 ( .A(n342), .ZN(n93) );
  OAI211_X1 U237 ( .C1(Rst), .C2(n349), .A(n319), .B(n313), .ZN(N175) );
  AND2_X1 U238 ( .A1(n356), .A2(n351), .ZN(n350) );
  AND3_X1 U239 ( .A1(n351), .A2(n84), .A3(n95), .ZN(n364) );
  AND2_X1 U240 ( .A1(n346), .A2(n84), .ZN(N182) );
  INV_X1 U241 ( .A(n313), .ZN(n91) );
  NOR4_X1 U242 ( .A1(IR_IN[9]), .A2(IR_IN[8]), .A3(IR_IN[7]), .A4(IR_IN[6]), 
        .ZN(n339) );
  INV_X1 U243 ( .A(n315), .ZN(n85) );
  AOI221_X1 U244 ( .B1(n316), .B2(n84), .C1(Rst), .C2(ALUCODE[1]), .A(n317), 
        .ZN(n315) );
  OAI221_X1 U245 ( .B1(n89), .B2(n109), .C1(n327), .C2(n328), .A(n86), .ZN(
        n316) );
  NOR2_X1 U246 ( .A1(n112), .A2(IR_IN_31), .ZN(n340) );
  NOR2_X1 U247 ( .A1(IR_IN_26), .A2(IR_IN_27), .ZN(n341) );
  NOR3_X1 U248 ( .A1(n97), .A2(IR_IN_27), .A3(n94), .ZN(n356) );
  NOR2_X1 U249 ( .A1(n108), .A2(IR_IN[0]), .ZN(n324) );
  OAI221_X1 U250 ( .B1(Rst), .B2(n335), .C1(n193), .C2(n84), .A(n336), .ZN(
        n103) );
  OAI211_X1 U251 ( .C1(n337), .C2(n99), .A(n111), .B(n87), .ZN(n336) );
  AOI221_X1 U252 ( .B1(n340), .B2(n95), .C1(n96), .C2(n341), .A(n329), .ZN(
        n335) );
  AOI21_X1 U253 ( .B1(n325), .B2(n326), .A(n110), .ZN(n337) );
  NAND4_X1 U254 ( .A1(n342), .A2(n343), .A3(n344), .A4(n345), .ZN(n329) );
  AOI21_X1 U255 ( .B1(n346), .B2(IR_IN_26), .A(n347), .ZN(n345) );
  NAND4_X1 U256 ( .A1(IR_IN[2]), .A2(n324), .A3(n99), .A4(n348), .ZN(n344) );
  NOR4_X1 U257 ( .A1(IR_IN_30), .A2(n94), .A3(n109), .A4(n327), .ZN(n347) );
  NAND2_X1 U258 ( .A1(IR_IN_27), .A2(n97), .ZN(n327) );
  NOR2_X1 U259 ( .A1(IR_IN_29), .A2(IR_IN_31), .ZN(n355) );
  AOI22_X1 U260 ( .A1(n323), .A2(IR_IN[0]), .B1(n324), .B2(n101), .ZN(n318) );
  INV_X1 U261 ( .A(n325), .ZN(n101) );
  AOI21_X1 U262 ( .B1(n322), .B2(n326), .A(IR_IN[1]), .ZN(n323) );
  INV_X1 U263 ( .A(IR_IN_28), .ZN(n94) );
  NAND2_X1 U264 ( .A1(IR_IN[3]), .A2(n338), .ZN(n326) );
  NAND2_X1 U265 ( .A1(n341), .A2(IR_IN_28), .ZN(n366) );
  OAI21_X1 U266 ( .B1(IR_IN_27), .B2(n97), .A(n366), .ZN(n367) );
  INV_X1 U267 ( .A(IR_IN_26), .ZN(n97) );
  OAI221_X1 U268 ( .B1(Rst), .B2(n330), .C1(n195), .C2(n84), .A(n331), .ZN(
        n105) );
  INV_X1 U269 ( .A(n326), .ZN(n100) );
  INV_X1 U270 ( .A(IR_IN[1]), .ZN(n108) );
  INV_X1 U271 ( .A(IR_IN_30), .ZN(n98) );
  INV_X1 U272 ( .A(IR_IN[2]), .ZN(n110) );
  AND4_X1 U273 ( .A1(n102), .A2(n106), .A3(IR_IN[5]), .A4(n339), .ZN(n338) );
  INV_X1 U274 ( .A(IR_IN[0]), .ZN(n111) );
  INV_X1 U275 ( .A(IR_IN_29), .ZN(n112) );
  OAI221_X1 U276 ( .B1(Rst), .B2(n332), .C1(n194), .C2(n84), .A(n333), .ZN(
        n104) );
  OR3_X1 U277 ( .A1(n319), .A2(n334), .A3(n322), .ZN(n333) );
  AOI21_X1 U278 ( .B1(n108), .B2(IR_IN[2]), .A(n324), .ZN(n334) );
  INV_X1 U279 ( .A(IR_IN[3]), .ZN(n107) );
  AND3_X1 U280 ( .A1(n94), .A2(n98), .A3(IR_IN_27), .ZN(n354) );
  INV_X1 U281 ( .A(IR_IN[4]), .ZN(n106) );
  INV_X1 U282 ( .A(IR_IN[10]), .ZN(n102) );
  NOR2_X1 U283 ( .A1(Rst), .A2(n358), .ZN(n277) );
  NOR2_X1 U284 ( .A1(Rst), .A2(n359), .ZN(n278) );
  NOR2_X1 U285 ( .A1(Rst), .A2(n360), .ZN(n279) );
  NOR2_X1 U286 ( .A1(Rst), .A2(n361), .ZN(n280) );
  NOR2_X1 U287 ( .A1(Rst), .A2(n362), .ZN(n281) );
  NOR2_X1 U288 ( .A1(Rst), .A2(n276), .ZN(n282) );
  NOR2_X1 U289 ( .A1(Rst), .A2(n275), .ZN(n283) );
  INV_X1 U290 ( .A(Rst), .ZN(n84) );
  NAND2_X1 U291 ( .A1(N182), .A2(IR_IN_26), .ZN(n313) );
  NOR2_X1 U292 ( .A1(IR_IN_29), .A2(n314), .ZN(N176) );
  AND4_X1 U293 ( .A1(n330), .A2(n343), .A3(n332), .A4(n357), .ZN(n349) );
  AOI21_X1 U294 ( .B1(n93), .B2(n112), .A(n363), .ZN(n357) );
  AOI21_X1 U295 ( .B1(IR_IN_27), .B2(n327), .A(n328), .ZN(n363) );
endmodule


module Adder_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module Adder ( A, B, reset, Cin, O, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  input reset, Cin;
  output Cout;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61,
         N62, N63, N64, N65, n17, n18, n19, n20;
  assign Cout = O[31];

  Adder_DW01_add_0 add_1_root_add_26_2 ( .A(A), .B(B), .CI(Cin), .SUM({N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, 
        N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, 
        N36, N35, N34}) );
  BUF_X1 U2 ( .A(n20), .Z(n17) );
  BUF_X1 U3 ( .A(n20), .Z(n18) );
  BUF_X1 U4 ( .A(n20), .Z(n19) );
  INV_X1 U5 ( .A(reset), .ZN(n20) );
  AND2_X1 U6 ( .A1(N34), .A2(n17), .ZN(O[0]) );
  AND2_X1 U7 ( .A1(N35), .A2(n17), .ZN(O[1]) );
  AND2_X1 U8 ( .A1(N36), .A2(n18), .ZN(O[2]) );
  AND2_X1 U9 ( .A1(N44), .A2(n17), .ZN(O[10]) );
  AND2_X1 U10 ( .A1(N45), .A2(n17), .ZN(O[11]) );
  AND2_X1 U11 ( .A1(N46), .A2(n17), .ZN(O[12]) );
  AND2_X1 U12 ( .A1(N47), .A2(n17), .ZN(O[13]) );
  AND2_X1 U13 ( .A1(N48), .A2(n17), .ZN(O[14]) );
  AND2_X1 U14 ( .A1(N49), .A2(n17), .ZN(O[15]) );
  AND2_X1 U15 ( .A1(N50), .A2(n17), .ZN(O[16]) );
  AND2_X1 U16 ( .A1(N51), .A2(n17), .ZN(O[17]) );
  AND2_X1 U17 ( .A1(N52), .A2(n17), .ZN(O[18]) );
  AND2_X1 U18 ( .A1(N53), .A2(n17), .ZN(O[19]) );
  AND2_X1 U19 ( .A1(N54), .A2(n18), .ZN(O[20]) );
  AND2_X1 U20 ( .A1(N55), .A2(n18), .ZN(O[21]) );
  AND2_X1 U21 ( .A1(N56), .A2(n18), .ZN(O[22]) );
  AND2_X1 U22 ( .A1(N57), .A2(n18), .ZN(O[23]) );
  AND2_X1 U23 ( .A1(N58), .A2(n18), .ZN(O[24]) );
  AND2_X1 U24 ( .A1(N59), .A2(n18), .ZN(O[25]) );
  AND2_X1 U25 ( .A1(N60), .A2(n18), .ZN(O[26]) );
  AND2_X1 U26 ( .A1(N61), .A2(n18), .ZN(O[27]) );
  AND2_X1 U27 ( .A1(N62), .A2(n18), .ZN(O[28]) );
  AND2_X1 U28 ( .A1(N63), .A2(n18), .ZN(O[29]) );
  AND2_X1 U29 ( .A1(N64), .A2(n18), .ZN(O[30]) );
  AND2_X1 U30 ( .A1(N37), .A2(n19), .ZN(O[3]) );
  AND2_X1 U31 ( .A1(N38), .A2(n19), .ZN(O[4]) );
  AND2_X1 U32 ( .A1(N39), .A2(n19), .ZN(O[5]) );
  AND2_X1 U33 ( .A1(N40), .A2(n19), .ZN(O[6]) );
  AND2_X1 U34 ( .A1(N41), .A2(n19), .ZN(O[7]) );
  AND2_X1 U35 ( .A1(N42), .A2(n19), .ZN(O[8]) );
  AND2_X1 U36 ( .A1(N43), .A2(n19), .ZN(O[9]) );
  AND2_X1 U37 ( .A1(N65), .A2(n19), .ZN(O[31]) );
endmodule


module IR ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n31, n32, n33, n34, n35, n97, n98, n99, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344;

  DFF_X1 \temp_reg[28]  ( .D(n66), .CK(clock), .Q(o[28]), .QN(n98) );
  DFF_X1 \temp_reg[23]  ( .D(n73), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[21]  ( .D(n75), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[25]  ( .D(n71), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[26]  ( .D(n65), .CK(clock), .Q(o[26]), .QN(n99) );
  DFF_X1 \temp_reg[30]  ( .D(n67), .CK(clock), .Q(o[30]), .QN(n97) );
  DFF_X1 \temp_reg[24]  ( .D(n72), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[5]  ( .D(n91), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[7]  ( .D(n89), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[8]  ( .D(n88), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[9]  ( .D(n87), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[10]  ( .D(n86), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[4]  ( .D(n92), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[11]  ( .D(n85), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[13]  ( .D(n83), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[14]  ( .D(n82), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[12]  ( .D(n84), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[6]  ( .D(n90), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[3]  ( .D(n93), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[1]  ( .D(n95), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n64) );
  DFF_X1 \temp_reg[2]  ( .D(n94), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[0]  ( .D(n96), .CK(clock), .Q(o[0]), .QN(n36) );
  DFF_X1 \temp_reg[20]  ( .D(n76), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n77), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[27]  ( .D(n70), .CK(clock), .Q(o[27]), .QN(n62) );
  DFF_X1 \temp_reg[29]  ( .D(n69), .CK(clock), .Q(o[29]), .QN(n63) );
  DFF_X1 \temp_reg[18]  ( .D(n78), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[16]  ( .D(n80), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[17]  ( .D(n79), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[15]  ( .D(n81), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[22]  ( .D(n74), .CK(clock), .Q(o[22]), .QN(n58) );
  INV_X1 U3 ( .A(reset), .ZN(n315) );
  BUF_X2 U4 ( .A(n32), .Z(n309) );
  BUF_X1 U5 ( .A(n32), .Z(n311) );
  BUF_X1 U6 ( .A(n31), .Z(n313) );
  BUF_X1 U7 ( .A(n31), .Z(n312) );
  BUF_X1 U8 ( .A(n31), .Z(n314) );
  INV_X1 U9 ( .A(i[15]), .ZN(n329) );
  INV_X1 U10 ( .A(i[18]), .ZN(n326) );
  INV_X1 U11 ( .A(i[19]), .ZN(n325) );
  INV_X1 U12 ( .A(i[20]), .ZN(n324) );
  INV_X1 U13 ( .A(i[21]), .ZN(n323) );
  INV_X1 U14 ( .A(i[23]), .ZN(n321) );
  INV_X1 U15 ( .A(i[0]), .ZN(n344) );
  INV_X1 U16 ( .A(i[2]), .ZN(n342) );
  INV_X1 U17 ( .A(i[1]), .ZN(n343) );
  INV_X1 U18 ( .A(i[3]), .ZN(n341) );
  INV_X1 U19 ( .A(i[6]), .ZN(n338) );
  INV_X1 U20 ( .A(i[11]), .ZN(n333) );
  INV_X1 U21 ( .A(i[4]), .ZN(n340) );
  INV_X1 U22 ( .A(i[10]), .ZN(n334) );
  INV_X1 U23 ( .A(i[9]), .ZN(n335) );
  INV_X1 U24 ( .A(i[8]), .ZN(n336) );
  INV_X1 U25 ( .A(i[7]), .ZN(n337) );
  INV_X1 U26 ( .A(i[5]), .ZN(n339) );
  OAI22_X1 U27 ( .A1(n313), .A2(n53), .B1(n310), .B2(n327), .ZN(n79) );
  INV_X1 U28 ( .A(i[17]), .ZN(n327) );
  OAI22_X1 U29 ( .A1(n313), .A2(n52), .B1(n310), .B2(n328), .ZN(n80) );
  INV_X1 U30 ( .A(i[16]), .ZN(n328) );
  OAI22_X1 U31 ( .A1(n313), .A2(n48), .B1(n310), .B2(n332), .ZN(n84) );
  INV_X1 U32 ( .A(i[12]), .ZN(n332) );
  OAI22_X1 U33 ( .A1(n313), .A2(n50), .B1(n310), .B2(n330), .ZN(n82) );
  INV_X1 U34 ( .A(i[14]), .ZN(n330) );
  OAI22_X1 U35 ( .A1(n313), .A2(n49), .B1(n310), .B2(n331), .ZN(n83) );
  INV_X1 U36 ( .A(i[13]), .ZN(n331) );
  OAI22_X1 U37 ( .A1(n313), .A2(n58), .B1(n310), .B2(n322), .ZN(n74) );
  INV_X1 U38 ( .A(i[22]), .ZN(n322) );
  OAI22_X1 U39 ( .A1(n314), .A2(n63), .B1(n311), .B2(n317), .ZN(n69) );
  INV_X1 U40 ( .A(i[29]), .ZN(n317) );
  OAI22_X1 U41 ( .A1(n314), .A2(n62), .B1(n311), .B2(n318), .ZN(n70) );
  INV_X1 U42 ( .A(i[27]), .ZN(n318) );
  OAI22_X1 U43 ( .A1(n314), .A2(n64), .B1(n311), .B2(n316), .ZN(n68) );
  INV_X1 U44 ( .A(i[31]), .ZN(n316) );
  OAI22_X1 U45 ( .A1(n314), .A2(n60), .B1(n311), .B2(n320), .ZN(n72) );
  INV_X1 U46 ( .A(i[24]), .ZN(n320) );
  OAI22_X1 U47 ( .A1(n314), .A2(n61), .B1(n311), .B2(n319), .ZN(n71) );
  INV_X1 U48 ( .A(i[25]), .ZN(n319) );
  OAI211_X1 U49 ( .C1(n314), .C2(n97), .A(n315), .B(n33), .ZN(n67) );
  NAND2_X1 U50 ( .A1(i[30]), .A2(n312), .ZN(n33) );
  OAI211_X1 U51 ( .C1(n314), .C2(n99), .A(n315), .B(n35), .ZN(n65) );
  NAND2_X1 U52 ( .A1(i[26]), .A2(n312), .ZN(n35) );
  OAI211_X1 U53 ( .C1(n314), .C2(n98), .A(n315), .B(n34), .ZN(n66) );
  NAND2_X1 U54 ( .A1(i[28]), .A2(n312), .ZN(n34) );
  OR2_X1 U55 ( .A1(reset), .A2(load), .ZN(n31) );
  OAI22_X1 U56 ( .A1(n313), .A2(n36), .B1(n309), .B2(n344), .ZN(n96) );
  OAI22_X1 U57 ( .A1(n312), .A2(n37), .B1(n309), .B2(n343), .ZN(n95) );
  OAI22_X1 U58 ( .A1(n312), .A2(n38), .B1(n309), .B2(n342), .ZN(n94) );
  OAI22_X1 U59 ( .A1(n312), .A2(n39), .B1(n309), .B2(n341), .ZN(n93) );
  OAI22_X1 U60 ( .A1(n312), .A2(n40), .B1(n309), .B2(n340), .ZN(n92) );
  OAI22_X1 U61 ( .A1(n312), .A2(n41), .B1(n309), .B2(n339), .ZN(n91) );
  OAI22_X1 U62 ( .A1(n312), .A2(n42), .B1(n309), .B2(n338), .ZN(n90) );
  OAI22_X1 U63 ( .A1(n312), .A2(n43), .B1(n309), .B2(n337), .ZN(n89) );
  OAI22_X1 U64 ( .A1(n312), .A2(n44), .B1(n309), .B2(n336), .ZN(n88) );
  OAI22_X1 U65 ( .A1(n312), .A2(n45), .B1(n309), .B2(n335), .ZN(n87) );
  OAI22_X1 U66 ( .A1(n312), .A2(n46), .B1(n309), .B2(n334), .ZN(n86) );
  OAI22_X1 U67 ( .A1(n313), .A2(n47), .B1(n309), .B2(n333), .ZN(n85) );
  OAI22_X1 U68 ( .A1(n313), .A2(n51), .B1(n310), .B2(n329), .ZN(n81) );
  OAI22_X1 U69 ( .A1(n314), .A2(n59), .B1(n310), .B2(n321), .ZN(n73) );
  OAI22_X1 U70 ( .A1(n313), .A2(n57), .B1(n310), .B2(n323), .ZN(n75) );
  OAI22_X1 U71 ( .A1(n313), .A2(n56), .B1(n310), .B2(n324), .ZN(n76) );
  OAI22_X1 U72 ( .A1(n313), .A2(n55), .B1(n310), .B2(n325), .ZN(n77) );
  OAI22_X1 U73 ( .A1(n313), .A2(n54), .B1(n310), .B2(n326), .ZN(n78) );
  BUF_X2 U74 ( .A(n32), .Z(n310) );
  NAND2_X1 U75 ( .A1(load), .A2(n315), .ZN(n32) );
endmodule


module reg_12 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n329) );
  BUF_X1 U4 ( .A(n35), .Z(n328) );
  BUF_X1 U5 ( .A(n35), .Z(n330) );
  BUF_X1 U6 ( .A(n34), .Z(n331) );
  BUF_X1 U7 ( .A(n34), .Z(n332) );
  BUF_X1 U8 ( .A(n34), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n35) );
  OAI22_X1 U10 ( .A1(n333), .A2(n36), .B1(n330), .B2(n366), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n366) );
  OAI22_X1 U12 ( .A1(n333), .A2(n37), .B1(n330), .B2(n365), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n365) );
  OAI22_X1 U14 ( .A1(n333), .A2(n38), .B1(n330), .B2(n364), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n364) );
  OAI22_X1 U16 ( .A1(n333), .A2(n39), .B1(n330), .B2(n363), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n363) );
  OAI22_X1 U18 ( .A1(n333), .A2(n40), .B1(n330), .B2(n362), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n362) );
  OAI22_X1 U20 ( .A1(n333), .A2(n41), .B1(n330), .B2(n361), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n361) );
  OAI22_X1 U22 ( .A1(n333), .A2(n42), .B1(n330), .B2(n360), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n360) );
  OAI22_X1 U24 ( .A1(n332), .A2(n43), .B1(n330), .B2(n359), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n359) );
  OAI22_X1 U26 ( .A1(n332), .A2(n44), .B1(n329), .B2(n358), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n358) );
  OAI22_X1 U28 ( .A1(n332), .A2(n45), .B1(n329), .B2(n357), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n357) );
  OAI22_X1 U30 ( .A1(n332), .A2(n46), .B1(n329), .B2(n356), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n356) );
  OAI22_X1 U32 ( .A1(n332), .A2(n47), .B1(n329), .B2(n355), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n355) );
  OAI22_X1 U34 ( .A1(n332), .A2(n48), .B1(n329), .B2(n354), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n354) );
  OAI22_X1 U36 ( .A1(n332), .A2(n49), .B1(n329), .B2(n353), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n353) );
  OAI22_X1 U38 ( .A1(n332), .A2(n50), .B1(n329), .B2(n352), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n352) );
  OAI22_X1 U40 ( .A1(n332), .A2(n51), .B1(n329), .B2(n351), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n351) );
  OAI22_X1 U42 ( .A1(n332), .A2(n52), .B1(n329), .B2(n350), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n350) );
  OAI22_X1 U44 ( .A1(n332), .A2(n53), .B1(n329), .B2(n349), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n349) );
  OAI22_X1 U46 ( .A1(n332), .A2(n54), .B1(n329), .B2(n348), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n348) );
  OAI22_X1 U48 ( .A1(n332), .A2(n55), .B1(n329), .B2(n347), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n347) );
  OAI22_X1 U50 ( .A1(n331), .A2(n56), .B1(n328), .B2(n346), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n346) );
  OAI22_X1 U52 ( .A1(n331), .A2(n57), .B1(n328), .B2(n345), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n345) );
  OAI22_X1 U54 ( .A1(n331), .A2(n58), .B1(n328), .B2(n344), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n344) );
  OAI22_X1 U56 ( .A1(n331), .A2(n59), .B1(n328), .B2(n343), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n343) );
  OAI22_X1 U58 ( .A1(n331), .A2(n60), .B1(n328), .B2(n342), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n342) );
  OAI22_X1 U60 ( .A1(n331), .A2(n61), .B1(n328), .B2(n341), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n341) );
  OAI22_X1 U62 ( .A1(n331), .A2(n62), .B1(n328), .B2(n340), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n340) );
  OAI22_X1 U64 ( .A1(n331), .A2(n63), .B1(n328), .B2(n339), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n339) );
  OAI22_X1 U66 ( .A1(n331), .A2(n64), .B1(n328), .B2(n338), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n338) );
  OAI22_X1 U68 ( .A1(n331), .A2(n65), .B1(n328), .B2(n337), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n337) );
  OAI22_X1 U70 ( .A1(n331), .A2(n66), .B1(n328), .B2(n336), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n336) );
  OAI22_X1 U72 ( .A1(n331), .A2(n67), .B1(n328), .B2(n335), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n335) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n34) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module fetchUnit ( clock, reset, en1, BranchPC, BRANCHfromDECODE, Instruction, 
        PCtoIM, IRtoDecode, NPCtoDecode );
  input [31:0] BranchPC;
  input [31:0] Instruction;
  output [31:0] PCtoIM;
  output [31:0] IRtoDecode;
  output [31:0] NPCtoDecode;
  input clock, reset, en1, BRANCHfromDECODE;
  wire   LOAD, \MuxtoPc[9] , \MuxtoPc[8] , \MuxtoPc[7] , \MuxtoPc[6] ,
         \MuxtoPc[5] , \MuxtoPc[4] , \MuxtoPc[3] , \MuxtoPc[31] ,
         \MuxtoPc[30] , \MuxtoPc[2] , \MuxtoPc[29] , \MuxtoPc[28] ,
         \MuxtoPc[27] , \MuxtoPc[26] , \MuxtoPc[25] , \MuxtoPc[24] ,
         \MuxtoPc[23] , \MuxtoPc[22] , \MuxtoPc[21] , \MuxtoPc[20] ,
         \MuxtoPc[1] , \MuxtoPc[19] , \MuxtoPc[18] , \MuxtoPc[17] ,
         \MuxtoPc[16] , \MuxtoPc[15] , \MuxtoPc[14] , \MuxtoPc[13] ,
         \MuxtoPc[12] , \MuxtoPc[11] , \MuxtoPc[10] , \MuxtoPc[0] ;
  wire   [31:0] AddertoMux;

  Adder nxpc ( .A(PCtoIM), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .reset(reset), .Cin(1'b0), .O(AddertoMux) );
  Mux21_0 pcmux ( .a(BranchPC), .b(AddertoMux), .sel(BRANCHfromDECODE), .y({
        \MuxtoPc[31] , \MuxtoPc[30] , \MuxtoPc[29] , \MuxtoPc[28] , 
        \MuxtoPc[27] , \MuxtoPc[26] , \MuxtoPc[25] , \MuxtoPc[24] , 
        \MuxtoPc[23] , \MuxtoPc[22] , \MuxtoPc[21] , \MuxtoPc[20] , 
        \MuxtoPc[19] , \MuxtoPc[18] , \MuxtoPc[17] , \MuxtoPc[16] , 
        \MuxtoPc[15] , \MuxtoPc[14] , \MuxtoPc[13] , \MuxtoPc[12] , 
        \MuxtoPc[11] , \MuxtoPc[10] , \MuxtoPc[9] , \MuxtoPc[8] , \MuxtoPc[7] , 
        \MuxtoPc[6] , \MuxtoPc[5] , \MuxtoPc[4] , \MuxtoPc[3] , \MuxtoPc[2] , 
        \MuxtoPc[1] , \MuxtoPc[0] }) );
  IR InstrReg ( .clock(clock), .reset(LOAD), .load(en1), .i(Instruction), .o(
        IRtoDecode) );
  reg_0 PC ( .clock(clock), .reset(reset), .load(en1), .i({\MuxtoPc[31] , 
        \MuxtoPc[30] , \MuxtoPc[29] , \MuxtoPc[28] , \MuxtoPc[27] , 
        \MuxtoPc[26] , \MuxtoPc[25] , \MuxtoPc[24] , \MuxtoPc[23] , 
        \MuxtoPc[22] , \MuxtoPc[21] , \MuxtoPc[20] , \MuxtoPc[19] , 
        \MuxtoPc[18] , \MuxtoPc[17] , \MuxtoPc[16] , \MuxtoPc[15] , 
        \MuxtoPc[14] , \MuxtoPc[13] , \MuxtoPc[12] , \MuxtoPc[11] , 
        \MuxtoPc[10] , \MuxtoPc[9] , \MuxtoPc[8] , \MuxtoPc[7] , \MuxtoPc[6] , 
        \MuxtoPc[5] , \MuxtoPc[4] , \MuxtoPc[3] , \MuxtoPc[2] , \MuxtoPc[1] , 
        \MuxtoPc[0] }), .o(PCtoIM) );
  reg_12 NPC ( .clock(clock), .reset(reset), .load(en1), .i(AddertoMux), .o(
        NPCtoDecode) );
  OR2_X1 U2 ( .A1(BRANCHfromDECODE), .A2(reset), .ZN(LOAD) );
endmodule


module Mux41 ( a, b, c, d, sel, y );
  input [31:0] a;
  input [31:0] b;
  input [31:0] c;
  input [31:0] d;
  input [1:0] sel;
  output [31:0] y;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332;

  BUF_X1 U1 ( .A(n6), .Z(n323) );
  BUF_X1 U2 ( .A(n6), .Z(n324) );
  BUF_X1 U3 ( .A(n4), .Z(n329) );
  BUF_X1 U4 ( .A(n4), .Z(n330) );
  BUF_X1 U5 ( .A(n7), .Z(n320) );
  BUF_X1 U6 ( .A(n7), .Z(n321) );
  BUF_X1 U7 ( .A(n5), .Z(n326) );
  BUF_X1 U8 ( .A(n5), .Z(n327) );
  BUF_X1 U9 ( .A(n6), .Z(n325) );
  BUF_X1 U10 ( .A(n4), .Z(n331) );
  BUF_X1 U11 ( .A(n7), .Z(n322) );
  BUF_X1 U12 ( .A(n5), .Z(n328) );
  AOI22_X1 U13 ( .A1(a[3]), .A2(n325), .B1(b[3]), .B2(n322), .ZN(n18) );
  AOI22_X1 U14 ( .A1(a[4]), .A2(n325), .B1(b[4]), .B2(n322), .ZN(n16) );
  AOI22_X1 U15 ( .A1(a[0]), .A2(n323), .B1(b[0]), .B2(n320), .ZN(n68) );
  AOI22_X1 U16 ( .A1(a[1]), .A2(n323), .B1(b[1]), .B2(n320), .ZN(n46) );
  AOI22_X1 U17 ( .A1(a[2]), .A2(n324), .B1(b[2]), .B2(n321), .ZN(n24) );
  NAND2_X1 U18 ( .A1(n24), .A2(n25), .ZN(y[2]) );
  AOI22_X1 U19 ( .A1(c[2]), .A2(n330), .B1(d[2]), .B2(n327), .ZN(n25) );
  NAND2_X1 U20 ( .A1(n18), .A2(n19), .ZN(y[3]) );
  AOI22_X1 U21 ( .A1(c[3]), .A2(n331), .B1(d[3]), .B2(n328), .ZN(n19) );
  NAND2_X1 U22 ( .A1(n16), .A2(n17), .ZN(y[4]) );
  AOI22_X1 U23 ( .A1(c[4]), .A2(n331), .B1(d[4]), .B2(n328), .ZN(n17) );
  NAND2_X1 U24 ( .A1(n68), .A2(n69), .ZN(y[0]) );
  AOI22_X1 U25 ( .A1(c[0]), .A2(n329), .B1(d[0]), .B2(n326), .ZN(n69) );
  NAND2_X1 U26 ( .A1(n46), .A2(n47), .ZN(y[1]) );
  AOI22_X1 U27 ( .A1(c[1]), .A2(n329), .B1(d[1]), .B2(n326), .ZN(n47) );
  NAND2_X1 U28 ( .A1(n14), .A2(n15), .ZN(y[5]) );
  AOI22_X1 U29 ( .A1(a[5]), .A2(n325), .B1(b[5]), .B2(n322), .ZN(n14) );
  NAND2_X1 U30 ( .A1(n12), .A2(n13), .ZN(y[6]) );
  AOI22_X1 U31 ( .A1(a[6]), .A2(n325), .B1(b[6]), .B2(n322), .ZN(n12) );
  NAND2_X1 U32 ( .A1(n44), .A2(n45), .ZN(y[20]) );
  AOI22_X1 U33 ( .A1(a[20]), .A2(n324), .B1(b[20]), .B2(n321), .ZN(n44) );
  NAND2_X1 U34 ( .A1(n42), .A2(n43), .ZN(y[21]) );
  AOI22_X1 U35 ( .A1(a[21]), .A2(n324), .B1(b[21]), .B2(n321), .ZN(n42) );
  NAND2_X1 U36 ( .A1(n40), .A2(n41), .ZN(y[22]) );
  AOI22_X1 U37 ( .A1(a[22]), .A2(n324), .B1(b[22]), .B2(n321), .ZN(n40) );
  NAND2_X1 U38 ( .A1(n38), .A2(n39), .ZN(y[23]) );
  AOI22_X1 U39 ( .A1(a[23]), .A2(n324), .B1(b[23]), .B2(n321), .ZN(n38) );
  NAND2_X1 U40 ( .A1(n36), .A2(n37), .ZN(y[24]) );
  AOI22_X1 U41 ( .A1(a[24]), .A2(n324), .B1(b[24]), .B2(n321), .ZN(n36) );
  NAND2_X1 U42 ( .A1(n34), .A2(n35), .ZN(y[25]) );
  AOI22_X1 U43 ( .A1(a[25]), .A2(n324), .B1(b[25]), .B2(n321), .ZN(n34) );
  NAND2_X1 U44 ( .A1(n32), .A2(n33), .ZN(y[26]) );
  AOI22_X1 U45 ( .A1(a[26]), .A2(n324), .B1(b[26]), .B2(n321), .ZN(n32) );
  NAND2_X1 U46 ( .A1(n30), .A2(n31), .ZN(y[27]) );
  AOI22_X1 U47 ( .A1(a[27]), .A2(n324), .B1(b[27]), .B2(n321), .ZN(n30) );
  NAND2_X1 U48 ( .A1(n28), .A2(n29), .ZN(y[28]) );
  AOI22_X1 U49 ( .A1(a[28]), .A2(n324), .B1(b[28]), .B2(n321), .ZN(n28) );
  NAND2_X1 U50 ( .A1(n26), .A2(n27), .ZN(y[29]) );
  AOI22_X1 U51 ( .A1(a[29]), .A2(n324), .B1(b[29]), .B2(n321), .ZN(n26) );
  NAND2_X1 U52 ( .A1(n22), .A2(n23), .ZN(y[30]) );
  AOI22_X1 U53 ( .A1(a[30]), .A2(n324), .B1(b[30]), .B2(n321), .ZN(n22) );
  NAND2_X1 U54 ( .A1(n20), .A2(n21), .ZN(y[31]) );
  AOI22_X1 U55 ( .A1(a[31]), .A2(n325), .B1(b[31]), .B2(n322), .ZN(n20) );
  NAND2_X1 U56 ( .A1(n10), .A2(n11), .ZN(y[7]) );
  AOI22_X1 U57 ( .A1(a[7]), .A2(n325), .B1(b[7]), .B2(n322), .ZN(n10) );
  NAND2_X1 U58 ( .A1(n8), .A2(n9), .ZN(y[8]) );
  AOI22_X1 U59 ( .A1(a[8]), .A2(n325), .B1(b[8]), .B2(n322), .ZN(n8) );
  NAND2_X1 U60 ( .A1(n2), .A2(n3), .ZN(y[9]) );
  AOI22_X1 U61 ( .A1(a[9]), .A2(n325), .B1(b[9]), .B2(n322), .ZN(n2) );
  NAND2_X1 U62 ( .A1(n66), .A2(n67), .ZN(y[10]) );
  AOI22_X1 U63 ( .A1(a[10]), .A2(n323), .B1(b[10]), .B2(n320), .ZN(n66) );
  NAND2_X1 U64 ( .A1(n64), .A2(n65), .ZN(y[11]) );
  AOI22_X1 U65 ( .A1(a[11]), .A2(n323), .B1(b[11]), .B2(n320), .ZN(n64) );
  NAND2_X1 U66 ( .A1(n62), .A2(n63), .ZN(y[12]) );
  AOI22_X1 U67 ( .A1(a[12]), .A2(n323), .B1(b[12]), .B2(n320), .ZN(n62) );
  NAND2_X1 U68 ( .A1(n60), .A2(n61), .ZN(y[13]) );
  AOI22_X1 U69 ( .A1(a[13]), .A2(n323), .B1(b[13]), .B2(n320), .ZN(n60) );
  NAND2_X1 U70 ( .A1(n58), .A2(n59), .ZN(y[14]) );
  AOI22_X1 U71 ( .A1(a[14]), .A2(n323), .B1(b[14]), .B2(n320), .ZN(n58) );
  NAND2_X1 U72 ( .A1(n56), .A2(n57), .ZN(y[15]) );
  AOI22_X1 U73 ( .A1(a[15]), .A2(n323), .B1(b[15]), .B2(n320), .ZN(n56) );
  NAND2_X1 U74 ( .A1(n54), .A2(n55), .ZN(y[16]) );
  AOI22_X1 U75 ( .A1(a[16]), .A2(n323), .B1(b[16]), .B2(n320), .ZN(n54) );
  NAND2_X1 U76 ( .A1(n52), .A2(n53), .ZN(y[17]) );
  AOI22_X1 U77 ( .A1(a[17]), .A2(n323), .B1(b[17]), .B2(n320), .ZN(n52) );
  NAND2_X1 U78 ( .A1(n50), .A2(n51), .ZN(y[18]) );
  AOI22_X1 U79 ( .A1(a[18]), .A2(n323), .B1(b[18]), .B2(n320), .ZN(n50) );
  NAND2_X1 U80 ( .A1(n48), .A2(n49), .ZN(y[19]) );
  AOI22_X1 U81 ( .A1(a[19]), .A2(n323), .B1(b[19]), .B2(n320), .ZN(n48) );
  NOR2_X1 U82 ( .A1(sel[0]), .A2(sel[1]), .ZN(n6) );
  NOR2_X1 U83 ( .A1(n332), .A2(sel[1]), .ZN(n7) );
  AND2_X1 U84 ( .A1(sel[1]), .A2(n332), .ZN(n4) );
  AND2_X1 U85 ( .A1(sel[0]), .A2(sel[1]), .ZN(n5) );
  INV_X1 U86 ( .A(sel[0]), .ZN(n332) );
  AOI22_X1 U87 ( .A1(c[5]), .A2(n331), .B1(d[5]), .B2(n328), .ZN(n15) );
  AOI22_X1 U88 ( .A1(c[6]), .A2(n331), .B1(d[6]), .B2(n328), .ZN(n13) );
  AOI22_X1 U89 ( .A1(c[7]), .A2(n331), .B1(d[7]), .B2(n328), .ZN(n11) );
  AOI22_X1 U90 ( .A1(c[8]), .A2(n331), .B1(d[8]), .B2(n328), .ZN(n9) );
  AOI22_X1 U91 ( .A1(c[9]), .A2(n331), .B1(d[9]), .B2(n328), .ZN(n3) );
  AOI22_X1 U92 ( .A1(c[10]), .A2(n329), .B1(d[10]), .B2(n326), .ZN(n67) );
  AOI22_X1 U93 ( .A1(c[11]), .A2(n329), .B1(d[11]), .B2(n326), .ZN(n65) );
  AOI22_X1 U94 ( .A1(c[12]), .A2(n329), .B1(d[12]), .B2(n326), .ZN(n63) );
  AOI22_X1 U95 ( .A1(c[13]), .A2(n329), .B1(d[13]), .B2(n326), .ZN(n61) );
  AOI22_X1 U96 ( .A1(c[14]), .A2(n329), .B1(d[14]), .B2(n326), .ZN(n59) );
  AOI22_X1 U97 ( .A1(c[15]), .A2(n329), .B1(d[15]), .B2(n326), .ZN(n57) );
  AOI22_X1 U98 ( .A1(c[16]), .A2(n329), .B1(d[16]), .B2(n326), .ZN(n55) );
  AOI22_X1 U99 ( .A1(c[17]), .A2(n329), .B1(d[17]), .B2(n326), .ZN(n53) );
  AOI22_X1 U100 ( .A1(c[18]), .A2(n329), .B1(d[18]), .B2(n326), .ZN(n51) );
  AOI22_X1 U101 ( .A1(c[19]), .A2(n329), .B1(d[19]), .B2(n326), .ZN(n49) );
  AOI22_X1 U102 ( .A1(c[20]), .A2(n330), .B1(d[20]), .B2(n327), .ZN(n45) );
  AOI22_X1 U103 ( .A1(c[21]), .A2(n330), .B1(d[21]), .B2(n327), .ZN(n43) );
  AOI22_X1 U104 ( .A1(c[22]), .A2(n330), .B1(d[22]), .B2(n327), .ZN(n41) );
  AOI22_X1 U105 ( .A1(c[23]), .A2(n330), .B1(d[23]), .B2(n327), .ZN(n39) );
  AOI22_X1 U106 ( .A1(c[24]), .A2(n330), .B1(d[24]), .B2(n327), .ZN(n37) );
  AOI22_X1 U107 ( .A1(c[25]), .A2(n330), .B1(d[25]), .B2(n327), .ZN(n35) );
  AOI22_X1 U108 ( .A1(c[26]), .A2(n330), .B1(d[26]), .B2(n327), .ZN(n33) );
  AOI22_X1 U109 ( .A1(c[27]), .A2(n330), .B1(d[27]), .B2(n327), .ZN(n31) );
  AOI22_X1 U110 ( .A1(c[28]), .A2(n330), .B1(d[28]), .B2(n327), .ZN(n29) );
  AOI22_X1 U111 ( .A1(c[29]), .A2(n330), .B1(d[29]), .B2(n327), .ZN(n27) );
  AOI22_X1 U112 ( .A1(c[30]), .A2(n330), .B1(d[30]), .B2(n327), .ZN(n23) );
  AOI22_X1 U113 ( .A1(c[31]), .A2(n331), .B1(d[31]), .B2(n328), .ZN(n21) );
endmodule


module BranchUnit ( a, sel, y );
  input [31:0] a;
  input sel;
  output y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NOR4_X1 U2 ( .A1(a[9]), .A2(a[8]), .A3(a[7]), .A4(a[6]), .ZN(n11) );
  NOR4_X1 U3 ( .A1(a[27]), .A2(a[26]), .A3(a[25]), .A4(a[24]), .ZN(n8) );
  NOR4_X1 U4 ( .A1(a[30]), .A2(a[2]), .A3(a[29]), .A4(a[28]), .ZN(n9) );
  NOR4_X1 U5 ( .A1(a[5]), .A2(a[4]), .A3(a[3]), .A4(a[31]), .ZN(n10) );
  NOR4_X1 U6 ( .A1(a[12]), .A2(a[11]), .A3(a[10]), .A4(a[0]), .ZN(n4) );
  NOR4_X1 U7 ( .A1(a[23]), .A2(a[22]), .A3(a[21]), .A4(a[20]), .ZN(n7) );
  NOR4_X1 U8 ( .A1(a[16]), .A2(a[15]), .A3(a[14]), .A4(a[13]), .ZN(n5) );
  NOR4_X1 U9 ( .A1(a[1]), .A2(a[19]), .A3(a[18]), .A4(a[17]), .ZN(n6) );
  NAND4_X1 U10 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(n3) );
  NOR2_X1 U11 ( .A1(n2), .A2(n3), .ZN(n1) );
  NAND4_X1 U12 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n2) );
  XNOR2_X1 U13 ( .A(sel), .B(n1), .ZN(y) );
endmodule


module reg_11 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n367), .Z(n329) );
  BUF_X1 U4 ( .A(n367), .Z(n328) );
  BUF_X1 U5 ( .A(n367), .Z(n330) );
  BUF_X1 U6 ( .A(n368), .Z(n331) );
  BUF_X1 U7 ( .A(n368), .Z(n332) );
  BUF_X1 U8 ( .A(n368), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n367) );
  OAI22_X1 U10 ( .A1(n333), .A2(n36), .B1(n330), .B2(n335), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n335) );
  OAI22_X1 U12 ( .A1(n333), .A2(n37), .B1(n330), .B2(n336), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n336) );
  OAI22_X1 U14 ( .A1(n333), .A2(n38), .B1(n330), .B2(n337), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n337) );
  OAI22_X1 U16 ( .A1(n333), .A2(n39), .B1(n330), .B2(n338), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n338) );
  OAI22_X1 U18 ( .A1(n333), .A2(n40), .B1(n330), .B2(n339), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n339) );
  OAI22_X1 U20 ( .A1(n333), .A2(n41), .B1(n330), .B2(n340), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n340) );
  OAI22_X1 U22 ( .A1(n333), .A2(n42), .B1(n330), .B2(n341), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n341) );
  OAI22_X1 U24 ( .A1(n332), .A2(n43), .B1(n330), .B2(n342), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n342) );
  OAI22_X1 U26 ( .A1(n332), .A2(n44), .B1(n329), .B2(n343), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n343) );
  OAI22_X1 U28 ( .A1(n332), .A2(n45), .B1(n329), .B2(n344), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n344) );
  OAI22_X1 U30 ( .A1(n332), .A2(n46), .B1(n329), .B2(n345), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n345) );
  OAI22_X1 U32 ( .A1(n332), .A2(n47), .B1(n329), .B2(n346), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n346) );
  OAI22_X1 U34 ( .A1(n332), .A2(n48), .B1(n329), .B2(n347), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n347) );
  OAI22_X1 U36 ( .A1(n332), .A2(n49), .B1(n329), .B2(n348), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n348) );
  OAI22_X1 U38 ( .A1(n332), .A2(n50), .B1(n329), .B2(n349), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n349) );
  OAI22_X1 U40 ( .A1(n332), .A2(n51), .B1(n329), .B2(n350), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n350) );
  OAI22_X1 U42 ( .A1(n332), .A2(n52), .B1(n329), .B2(n351), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n351) );
  OAI22_X1 U44 ( .A1(n332), .A2(n53), .B1(n329), .B2(n352), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n352) );
  OAI22_X1 U46 ( .A1(n332), .A2(n54), .B1(n329), .B2(n353), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n353) );
  OAI22_X1 U48 ( .A1(n332), .A2(n55), .B1(n329), .B2(n354), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n354) );
  OAI22_X1 U50 ( .A1(n331), .A2(n56), .B1(n328), .B2(n355), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n355) );
  OAI22_X1 U52 ( .A1(n331), .A2(n57), .B1(n328), .B2(n356), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n356) );
  OAI22_X1 U54 ( .A1(n331), .A2(n58), .B1(n328), .B2(n357), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n357) );
  OAI22_X1 U56 ( .A1(n331), .A2(n59), .B1(n328), .B2(n358), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n358) );
  OAI22_X1 U58 ( .A1(n331), .A2(n60), .B1(n328), .B2(n359), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n359) );
  OAI22_X1 U60 ( .A1(n331), .A2(n61), .B1(n328), .B2(n360), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n360) );
  OAI22_X1 U62 ( .A1(n331), .A2(n62), .B1(n328), .B2(n361), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n361) );
  OAI22_X1 U64 ( .A1(n331), .A2(n63), .B1(n328), .B2(n362), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n362) );
  OAI22_X1 U66 ( .A1(n331), .A2(n64), .B1(n328), .B2(n363), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n363) );
  OAI22_X1 U68 ( .A1(n331), .A2(n65), .B1(n328), .B2(n364), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n364) );
  OAI22_X1 U70 ( .A1(n331), .A2(n66), .B1(n328), .B2(n365), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n365) );
  OAI22_X1 U72 ( .A1(n331), .A2(n67), .B1(n328), .B2(n366), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n366) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n368) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module reg_10 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n327) );
  BUF_X1 U4 ( .A(n35), .Z(n326) );
  BUF_X1 U5 ( .A(n35), .Z(n328) );
  BUF_X1 U6 ( .A(n34), .Z(n329) );
  BUF_X1 U7 ( .A(n34), .Z(n330) );
  BUF_X1 U8 ( .A(n34), .Z(n331) );
  NAND2_X1 U9 ( .A1(n332), .A2(n329), .ZN(n35) );
  OAI22_X1 U10 ( .A1(n330), .A2(n44), .B1(n327), .B2(n364), .ZN(n91) );
  INV_X1 U11 ( .A(i[8]), .ZN(n364) );
  OAI22_X1 U12 ( .A1(n330), .A2(n47), .B1(n327), .B2(n361), .ZN(n88) );
  INV_X1 U13 ( .A(i[11]), .ZN(n361) );
  OAI22_X1 U14 ( .A1(n330), .A2(n49), .B1(n327), .B2(n359), .ZN(n86) );
  INV_X1 U15 ( .A(i[13]), .ZN(n359) );
  OAI22_X1 U16 ( .A1(n330), .A2(n51), .B1(n327), .B2(n357), .ZN(n84) );
  INV_X1 U17 ( .A(i[15]), .ZN(n357) );
  OAI22_X1 U18 ( .A1(n330), .A2(n53), .B1(n327), .B2(n355), .ZN(n82) );
  INV_X1 U19 ( .A(i[17]), .ZN(n355) );
  OAI22_X1 U20 ( .A1(n330), .A2(n55), .B1(n327), .B2(n353), .ZN(n80) );
  INV_X1 U21 ( .A(i[19]), .ZN(n353) );
  OAI22_X1 U22 ( .A1(n329), .A2(n56), .B1(n326), .B2(n352), .ZN(n79) );
  INV_X1 U23 ( .A(i[20]), .ZN(n352) );
  OAI22_X1 U24 ( .A1(n329), .A2(n58), .B1(n326), .B2(n350), .ZN(n77) );
  INV_X1 U25 ( .A(i[22]), .ZN(n350) );
  OAI22_X1 U26 ( .A1(n329), .A2(n63), .B1(n326), .B2(n345), .ZN(n72) );
  INV_X1 U27 ( .A(i[27]), .ZN(n345) );
  OAI22_X1 U28 ( .A1(n329), .A2(n66), .B1(n326), .B2(n342), .ZN(n69) );
  INV_X1 U29 ( .A(i[30]), .ZN(n342) );
  OAI22_X1 U30 ( .A1(n331), .A2(n36), .B1(n328), .B2(n340), .ZN(n99) );
  INV_X1 U31 ( .A(i[0]), .ZN(n340) );
  OAI22_X1 U32 ( .A1(n331), .A2(n42), .B1(n328), .B2(n334), .ZN(n93) );
  INV_X1 U33 ( .A(i[6]), .ZN(n334) );
  OAI22_X1 U34 ( .A1(n329), .A2(n60), .B1(n326), .B2(n348), .ZN(n75) );
  INV_X1 U35 ( .A(i[24]), .ZN(n348) );
  OAI22_X1 U36 ( .A1(n329), .A2(n64), .B1(n326), .B2(n344), .ZN(n71) );
  INV_X1 U37 ( .A(i[28]), .ZN(n344) );
  OAI22_X1 U38 ( .A1(n329), .A2(n67), .B1(n326), .B2(n341), .ZN(n68) );
  INV_X1 U39 ( .A(i[31]), .ZN(n341) );
  OAI22_X1 U40 ( .A1(n331), .A2(n39), .B1(n328), .B2(n337), .ZN(n96) );
  INV_X1 U41 ( .A(i[3]), .ZN(n337) );
  OAI22_X1 U42 ( .A1(n330), .A2(n43), .B1(n328), .B2(n333), .ZN(n92) );
  INV_X1 U43 ( .A(i[7]), .ZN(n333) );
  OAI22_X1 U44 ( .A1(n330), .A2(n46), .B1(n327), .B2(n362), .ZN(n89) );
  INV_X1 U45 ( .A(i[10]), .ZN(n362) );
  OAI22_X1 U46 ( .A1(n330), .A2(n50), .B1(n327), .B2(n358), .ZN(n85) );
  INV_X1 U47 ( .A(i[14]), .ZN(n358) );
  OAI22_X1 U48 ( .A1(n330), .A2(n54), .B1(n327), .B2(n354), .ZN(n81) );
  INV_X1 U49 ( .A(i[18]), .ZN(n354) );
  OAI22_X1 U50 ( .A1(n329), .A2(n57), .B1(n326), .B2(n351), .ZN(n78) );
  INV_X1 U51 ( .A(i[21]), .ZN(n351) );
  OAI22_X1 U52 ( .A1(n329), .A2(n61), .B1(n326), .B2(n347), .ZN(n74) );
  INV_X1 U53 ( .A(i[25]), .ZN(n347) );
  OAI22_X1 U54 ( .A1(n329), .A2(n65), .B1(n326), .B2(n343), .ZN(n70) );
  INV_X1 U55 ( .A(i[29]), .ZN(n343) );
  OAI22_X1 U56 ( .A1(n331), .A2(n38), .B1(n328), .B2(n338), .ZN(n97) );
  INV_X1 U57 ( .A(i[2]), .ZN(n338) );
  OAI22_X1 U58 ( .A1(n331), .A2(n40), .B1(n328), .B2(n336), .ZN(n95) );
  INV_X1 U59 ( .A(i[4]), .ZN(n336) );
  OAI22_X1 U60 ( .A1(n329), .A2(n62), .B1(n326), .B2(n346), .ZN(n73) );
  INV_X1 U61 ( .A(i[26]), .ZN(n346) );
  OAI22_X1 U62 ( .A1(n331), .A2(n37), .B1(n328), .B2(n339), .ZN(n98) );
  INV_X1 U63 ( .A(i[1]), .ZN(n339) );
  OAI22_X1 U64 ( .A1(n331), .A2(n41), .B1(n328), .B2(n335), .ZN(n94) );
  INV_X1 U65 ( .A(i[5]), .ZN(n335) );
  OAI22_X1 U66 ( .A1(n330), .A2(n45), .B1(n327), .B2(n363), .ZN(n90) );
  INV_X1 U67 ( .A(i[9]), .ZN(n363) );
  OAI22_X1 U68 ( .A1(n330), .A2(n48), .B1(n327), .B2(n360), .ZN(n87) );
  INV_X1 U69 ( .A(i[12]), .ZN(n360) );
  OAI22_X1 U70 ( .A1(n330), .A2(n52), .B1(n327), .B2(n356), .ZN(n83) );
  INV_X1 U71 ( .A(i[16]), .ZN(n356) );
  OAI22_X1 U72 ( .A1(n329), .A2(n59), .B1(n326), .B2(n349), .ZN(n76) );
  INV_X1 U73 ( .A(i[23]), .ZN(n349) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n34) );
  INV_X1 U75 ( .A(reset), .ZN(n332) );
endmodule


module reg_9 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n367), .Z(n329) );
  BUF_X1 U4 ( .A(n367), .Z(n328) );
  BUF_X1 U5 ( .A(n367), .Z(n330) );
  BUF_X1 U6 ( .A(n368), .Z(n331) );
  BUF_X1 U7 ( .A(n368), .Z(n332) );
  BUF_X1 U8 ( .A(n368), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n367) );
  OAI22_X1 U10 ( .A1(n331), .A2(n60), .B1(n328), .B2(n350), .ZN(n75) );
  INV_X1 U11 ( .A(i[24]), .ZN(n350) );
  OAI22_X1 U12 ( .A1(n331), .A2(n61), .B1(n328), .B2(n349), .ZN(n74) );
  INV_X1 U13 ( .A(i[25]), .ZN(n349) );
  OAI22_X1 U14 ( .A1(n331), .A2(n62), .B1(n328), .B2(n348), .ZN(n73) );
  INV_X1 U15 ( .A(i[26]), .ZN(n348) );
  OAI22_X1 U16 ( .A1(n331), .A2(n63), .B1(n328), .B2(n347), .ZN(n72) );
  INV_X1 U17 ( .A(i[27]), .ZN(n347) );
  OAI22_X1 U18 ( .A1(n331), .A2(n64), .B1(n328), .B2(n346), .ZN(n71) );
  INV_X1 U19 ( .A(i[28]), .ZN(n346) );
  OAI22_X1 U20 ( .A1(n331), .A2(n65), .B1(n328), .B2(n345), .ZN(n70) );
  INV_X1 U21 ( .A(i[29]), .ZN(n345) );
  OAI22_X1 U22 ( .A1(n331), .A2(n66), .B1(n328), .B2(n344), .ZN(n69) );
  INV_X1 U23 ( .A(i[30]), .ZN(n344) );
  OAI22_X1 U24 ( .A1(n331), .A2(n67), .B1(n328), .B2(n343), .ZN(n68) );
  INV_X1 U25 ( .A(i[31]), .ZN(n343) );
  OAI22_X1 U26 ( .A1(n333), .A2(n36), .B1(n330), .B2(n342), .ZN(n99) );
  INV_X1 U27 ( .A(i[0]), .ZN(n342) );
  OAI22_X1 U28 ( .A1(n333), .A2(n37), .B1(n330), .B2(n341), .ZN(n98) );
  INV_X1 U29 ( .A(i[1]), .ZN(n341) );
  OAI22_X1 U30 ( .A1(n333), .A2(n38), .B1(n330), .B2(n340), .ZN(n97) );
  INV_X1 U31 ( .A(i[2]), .ZN(n340) );
  OAI22_X1 U32 ( .A1(n333), .A2(n39), .B1(n330), .B2(n339), .ZN(n96) );
  INV_X1 U33 ( .A(i[3]), .ZN(n339) );
  OAI22_X1 U34 ( .A1(n333), .A2(n40), .B1(n330), .B2(n338), .ZN(n95) );
  INV_X1 U35 ( .A(i[4]), .ZN(n338) );
  OAI22_X1 U36 ( .A1(n333), .A2(n41), .B1(n330), .B2(n337), .ZN(n94) );
  INV_X1 U37 ( .A(i[5]), .ZN(n337) );
  OAI22_X1 U38 ( .A1(n333), .A2(n42), .B1(n330), .B2(n336), .ZN(n93) );
  INV_X1 U39 ( .A(i[6]), .ZN(n336) );
  OAI22_X1 U40 ( .A1(n332), .A2(n43), .B1(n330), .B2(n335), .ZN(n92) );
  INV_X1 U41 ( .A(i[7]), .ZN(n335) );
  OAI22_X1 U42 ( .A1(n332), .A2(n44), .B1(n329), .B2(n366), .ZN(n91) );
  INV_X1 U43 ( .A(i[8]), .ZN(n366) );
  OAI22_X1 U44 ( .A1(n332), .A2(n45), .B1(n329), .B2(n365), .ZN(n90) );
  INV_X1 U45 ( .A(i[9]), .ZN(n365) );
  OAI22_X1 U46 ( .A1(n332), .A2(n46), .B1(n329), .B2(n364), .ZN(n89) );
  INV_X1 U47 ( .A(i[10]), .ZN(n364) );
  OAI22_X1 U48 ( .A1(n332), .A2(n47), .B1(n329), .B2(n363), .ZN(n88) );
  INV_X1 U49 ( .A(i[11]), .ZN(n363) );
  OAI22_X1 U50 ( .A1(n332), .A2(n48), .B1(n329), .B2(n362), .ZN(n87) );
  INV_X1 U51 ( .A(i[12]), .ZN(n362) );
  OAI22_X1 U52 ( .A1(n332), .A2(n49), .B1(n329), .B2(n361), .ZN(n86) );
  INV_X1 U53 ( .A(i[13]), .ZN(n361) );
  OAI22_X1 U54 ( .A1(n332), .A2(n50), .B1(n329), .B2(n360), .ZN(n85) );
  INV_X1 U55 ( .A(i[14]), .ZN(n360) );
  OAI22_X1 U56 ( .A1(n332), .A2(n51), .B1(n329), .B2(n359), .ZN(n84) );
  INV_X1 U57 ( .A(i[15]), .ZN(n359) );
  OAI22_X1 U58 ( .A1(n332), .A2(n52), .B1(n329), .B2(n358), .ZN(n83) );
  INV_X1 U59 ( .A(i[16]), .ZN(n358) );
  OAI22_X1 U60 ( .A1(n332), .A2(n53), .B1(n329), .B2(n357), .ZN(n82) );
  INV_X1 U61 ( .A(i[17]), .ZN(n357) );
  OAI22_X1 U62 ( .A1(n332), .A2(n54), .B1(n329), .B2(n356), .ZN(n81) );
  INV_X1 U63 ( .A(i[18]), .ZN(n356) );
  OAI22_X1 U64 ( .A1(n332), .A2(n55), .B1(n329), .B2(n355), .ZN(n80) );
  INV_X1 U65 ( .A(i[19]), .ZN(n355) );
  OAI22_X1 U66 ( .A1(n331), .A2(n56), .B1(n328), .B2(n354), .ZN(n79) );
  INV_X1 U67 ( .A(i[20]), .ZN(n354) );
  OAI22_X1 U68 ( .A1(n331), .A2(n57), .B1(n328), .B2(n353), .ZN(n78) );
  INV_X1 U69 ( .A(i[21]), .ZN(n353) );
  OAI22_X1 U70 ( .A1(n331), .A2(n58), .B1(n328), .B2(n352), .ZN(n77) );
  INV_X1 U71 ( .A(i[22]), .ZN(n352) );
  OAI22_X1 U72 ( .A1(n331), .A2(n59), .B1(n328), .B2(n351), .ZN(n76) );
  INV_X1 U73 ( .A(i[23]), .ZN(n351) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n368) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module reg_8 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n367), .Z(n329) );
  BUF_X1 U4 ( .A(n367), .Z(n328) );
  BUF_X1 U5 ( .A(n367), .Z(n330) );
  BUF_X1 U6 ( .A(n368), .Z(n331) );
  BUF_X1 U7 ( .A(n368), .Z(n332) );
  BUF_X1 U8 ( .A(n368), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n367) );
  OAI22_X1 U10 ( .A1(n333), .A2(n37), .B1(n330), .B2(n365), .ZN(n98) );
  INV_X1 U11 ( .A(i[1]), .ZN(n365) );
  OAI22_X1 U12 ( .A1(n333), .A2(n38), .B1(n330), .B2(n364), .ZN(n97) );
  INV_X1 U13 ( .A(i[2]), .ZN(n364) );
  OAI22_X1 U14 ( .A1(n333), .A2(n42), .B1(n330), .B2(n360), .ZN(n93) );
  INV_X1 U15 ( .A(i[6]), .ZN(n360) );
  OAI22_X1 U16 ( .A1(n332), .A2(n43), .B1(n330), .B2(n359), .ZN(n92) );
  INV_X1 U17 ( .A(i[7]), .ZN(n359) );
  OAI22_X1 U18 ( .A1(n332), .A2(n44), .B1(n329), .B2(n358), .ZN(n91) );
  INV_X1 U19 ( .A(i[8]), .ZN(n358) );
  OAI22_X1 U20 ( .A1(n332), .A2(n46), .B1(n329), .B2(n356), .ZN(n89) );
  INV_X1 U21 ( .A(i[10]), .ZN(n356) );
  OAI22_X1 U22 ( .A1(n332), .A2(n47), .B1(n329), .B2(n355), .ZN(n88) );
  INV_X1 U23 ( .A(i[11]), .ZN(n355) );
  OAI22_X1 U24 ( .A1(n332), .A2(n48), .B1(n329), .B2(n354), .ZN(n87) );
  INV_X1 U25 ( .A(i[12]), .ZN(n354) );
  OAI22_X1 U26 ( .A1(n332), .A2(n49), .B1(n329), .B2(n353), .ZN(n86) );
  INV_X1 U27 ( .A(i[13]), .ZN(n353) );
  OAI22_X1 U28 ( .A1(n332), .A2(n50), .B1(n329), .B2(n352), .ZN(n85) );
  INV_X1 U29 ( .A(i[14]), .ZN(n352) );
  OAI22_X1 U30 ( .A1(n332), .A2(n51), .B1(n329), .B2(n351), .ZN(n84) );
  INV_X1 U31 ( .A(i[15]), .ZN(n351) );
  OAI22_X1 U32 ( .A1(n332), .A2(n52), .B1(n329), .B2(n350), .ZN(n83) );
  INV_X1 U33 ( .A(i[16]), .ZN(n350) );
  OAI22_X1 U34 ( .A1(n332), .A2(n53), .B1(n329), .B2(n349), .ZN(n82) );
  INV_X1 U35 ( .A(i[17]), .ZN(n349) );
  OAI22_X1 U36 ( .A1(n332), .A2(n54), .B1(n329), .B2(n348), .ZN(n81) );
  INV_X1 U37 ( .A(i[18]), .ZN(n348) );
  OAI22_X1 U38 ( .A1(n332), .A2(n55), .B1(n329), .B2(n347), .ZN(n80) );
  INV_X1 U39 ( .A(i[19]), .ZN(n347) );
  OAI22_X1 U40 ( .A1(n331), .A2(n56), .B1(n328), .B2(n346), .ZN(n79) );
  INV_X1 U41 ( .A(i[20]), .ZN(n346) );
  OAI22_X1 U42 ( .A1(n331), .A2(n57), .B1(n328), .B2(n345), .ZN(n78) );
  INV_X1 U43 ( .A(i[21]), .ZN(n345) );
  OAI22_X1 U44 ( .A1(n331), .A2(n58), .B1(n328), .B2(n344), .ZN(n77) );
  INV_X1 U45 ( .A(i[22]), .ZN(n344) );
  OAI22_X1 U46 ( .A1(n331), .A2(n59), .B1(n328), .B2(n343), .ZN(n76) );
  INV_X1 U47 ( .A(i[23]), .ZN(n343) );
  OAI22_X1 U48 ( .A1(n331), .A2(n60), .B1(n328), .B2(n342), .ZN(n75) );
  INV_X1 U49 ( .A(i[24]), .ZN(n342) );
  OAI22_X1 U50 ( .A1(n331), .A2(n61), .B1(n328), .B2(n341), .ZN(n74) );
  INV_X1 U51 ( .A(i[25]), .ZN(n341) );
  OAI22_X1 U52 ( .A1(n331), .A2(n62), .B1(n328), .B2(n340), .ZN(n73) );
  INV_X1 U53 ( .A(i[26]), .ZN(n340) );
  OAI22_X1 U54 ( .A1(n331), .A2(n63), .B1(n328), .B2(n339), .ZN(n72) );
  INV_X1 U55 ( .A(i[27]), .ZN(n339) );
  OAI22_X1 U56 ( .A1(n331), .A2(n64), .B1(n328), .B2(n338), .ZN(n71) );
  INV_X1 U57 ( .A(i[28]), .ZN(n338) );
  OAI22_X1 U58 ( .A1(n331), .A2(n65), .B1(n328), .B2(n337), .ZN(n70) );
  INV_X1 U59 ( .A(i[29]), .ZN(n337) );
  OAI22_X1 U60 ( .A1(n331), .A2(n66), .B1(n328), .B2(n336), .ZN(n69) );
  INV_X1 U61 ( .A(i[30]), .ZN(n336) );
  OAI22_X1 U62 ( .A1(n331), .A2(n67), .B1(n328), .B2(n335), .ZN(n68) );
  INV_X1 U63 ( .A(i[31]), .ZN(n335) );
  OAI22_X1 U64 ( .A1(n333), .A2(n36), .B1(n330), .B2(n366), .ZN(n99) );
  INV_X1 U65 ( .A(i[0]), .ZN(n366) );
  OAI22_X1 U66 ( .A1(n333), .A2(n39), .B1(n330), .B2(n363), .ZN(n96) );
  INV_X1 U67 ( .A(i[3]), .ZN(n363) );
  OAI22_X1 U68 ( .A1(n333), .A2(n40), .B1(n330), .B2(n362), .ZN(n95) );
  INV_X1 U69 ( .A(i[4]), .ZN(n362) );
  OAI22_X1 U70 ( .A1(n333), .A2(n41), .B1(n330), .B2(n361), .ZN(n94) );
  INV_X1 U71 ( .A(i[5]), .ZN(n361) );
  OAI22_X1 U72 ( .A1(n332), .A2(n45), .B1(n329), .B2(n357), .ZN(n90) );
  INV_X1 U73 ( .A(i[9]), .ZN(n357) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n368) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module reg_7 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n367), .Z(n329) );
  BUF_X1 U4 ( .A(n367), .Z(n328) );
  BUF_X1 U5 ( .A(n367), .Z(n330) );
  BUF_X1 U6 ( .A(n368), .Z(n331) );
  BUF_X1 U7 ( .A(n368), .Z(n332) );
  BUF_X1 U8 ( .A(n368), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n367) );
  OAI22_X1 U10 ( .A1(n333), .A2(n38), .B1(n330), .B2(n336), .ZN(n97) );
  INV_X1 U11 ( .A(i[2]), .ZN(n336) );
  OAI22_X1 U12 ( .A1(n333), .A2(n39), .B1(n330), .B2(n337), .ZN(n96) );
  INV_X1 U13 ( .A(i[3]), .ZN(n337) );
  OAI22_X1 U14 ( .A1(n333), .A2(n40), .B1(n330), .B2(n339), .ZN(n95) );
  INV_X1 U15 ( .A(i[4]), .ZN(n339) );
  OAI22_X1 U16 ( .A1(n333), .A2(n36), .B1(n330), .B2(n335), .ZN(n99) );
  INV_X1 U17 ( .A(i[0]), .ZN(n335) );
  OAI22_X1 U18 ( .A1(n333), .A2(n37), .B1(n330), .B2(n338), .ZN(n98) );
  INV_X1 U19 ( .A(i[1]), .ZN(n338) );
  OAI22_X1 U20 ( .A1(n333), .A2(n41), .B1(n330), .B2(n340), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n340) );
  OAI22_X1 U22 ( .A1(n333), .A2(n42), .B1(n330), .B2(n341), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n341) );
  OAI22_X1 U24 ( .A1(n331), .A2(n56), .B1(n328), .B2(n355), .ZN(n79) );
  INV_X1 U25 ( .A(i[20]), .ZN(n355) );
  OAI22_X1 U26 ( .A1(n331), .A2(n57), .B1(n328), .B2(n356), .ZN(n78) );
  INV_X1 U27 ( .A(i[21]), .ZN(n356) );
  OAI22_X1 U28 ( .A1(n331), .A2(n58), .B1(n328), .B2(n357), .ZN(n77) );
  INV_X1 U29 ( .A(i[22]), .ZN(n357) );
  OAI22_X1 U30 ( .A1(n331), .A2(n59), .B1(n328), .B2(n358), .ZN(n76) );
  INV_X1 U31 ( .A(i[23]), .ZN(n358) );
  OAI22_X1 U32 ( .A1(n331), .A2(n60), .B1(n328), .B2(n359), .ZN(n75) );
  INV_X1 U33 ( .A(i[24]), .ZN(n359) );
  OAI22_X1 U34 ( .A1(n331), .A2(n61), .B1(n328), .B2(n360), .ZN(n74) );
  INV_X1 U35 ( .A(i[25]), .ZN(n360) );
  OAI22_X1 U36 ( .A1(n331), .A2(n62), .B1(n328), .B2(n361), .ZN(n73) );
  INV_X1 U37 ( .A(i[26]), .ZN(n361) );
  OAI22_X1 U38 ( .A1(n331), .A2(n63), .B1(n328), .B2(n362), .ZN(n72) );
  INV_X1 U39 ( .A(i[27]), .ZN(n362) );
  OAI22_X1 U40 ( .A1(n331), .A2(n64), .B1(n328), .B2(n363), .ZN(n71) );
  INV_X1 U41 ( .A(i[28]), .ZN(n363) );
  OAI22_X1 U42 ( .A1(n331), .A2(n65), .B1(n328), .B2(n364), .ZN(n70) );
  INV_X1 U43 ( .A(i[29]), .ZN(n364) );
  OAI22_X1 U44 ( .A1(n331), .A2(n66), .B1(n328), .B2(n365), .ZN(n69) );
  INV_X1 U45 ( .A(i[30]), .ZN(n365) );
  OAI22_X1 U46 ( .A1(n331), .A2(n67), .B1(n328), .B2(n366), .ZN(n68) );
  INV_X1 U47 ( .A(i[31]), .ZN(n366) );
  OAI22_X1 U48 ( .A1(n332), .A2(n43), .B1(n330), .B2(n342), .ZN(n92) );
  INV_X1 U49 ( .A(i[7]), .ZN(n342) );
  OAI22_X1 U50 ( .A1(n332), .A2(n44), .B1(n329), .B2(n343), .ZN(n91) );
  INV_X1 U51 ( .A(i[8]), .ZN(n343) );
  OAI22_X1 U52 ( .A1(n332), .A2(n45), .B1(n329), .B2(n344), .ZN(n90) );
  INV_X1 U53 ( .A(i[9]), .ZN(n344) );
  OAI22_X1 U54 ( .A1(n332), .A2(n46), .B1(n329), .B2(n345), .ZN(n89) );
  INV_X1 U55 ( .A(i[10]), .ZN(n345) );
  OAI22_X1 U56 ( .A1(n332), .A2(n47), .B1(n329), .B2(n346), .ZN(n88) );
  INV_X1 U57 ( .A(i[11]), .ZN(n346) );
  OAI22_X1 U58 ( .A1(n332), .A2(n48), .B1(n329), .B2(n347), .ZN(n87) );
  INV_X1 U59 ( .A(i[12]), .ZN(n347) );
  OAI22_X1 U60 ( .A1(n332), .A2(n49), .B1(n329), .B2(n348), .ZN(n86) );
  INV_X1 U61 ( .A(i[13]), .ZN(n348) );
  OAI22_X1 U62 ( .A1(n332), .A2(n50), .B1(n329), .B2(n349), .ZN(n85) );
  INV_X1 U63 ( .A(i[14]), .ZN(n349) );
  OAI22_X1 U64 ( .A1(n332), .A2(n51), .B1(n329), .B2(n350), .ZN(n84) );
  INV_X1 U65 ( .A(i[15]), .ZN(n350) );
  OAI22_X1 U66 ( .A1(n332), .A2(n52), .B1(n329), .B2(n351), .ZN(n83) );
  INV_X1 U67 ( .A(i[16]), .ZN(n351) );
  OAI22_X1 U68 ( .A1(n332), .A2(n53), .B1(n329), .B2(n352), .ZN(n82) );
  INV_X1 U69 ( .A(i[17]), .ZN(n352) );
  OAI22_X1 U70 ( .A1(n332), .A2(n54), .B1(n329), .B2(n353), .ZN(n81) );
  INV_X1 U71 ( .A(i[18]), .ZN(n353) );
  OAI22_X1 U72 ( .A1(n332), .A2(n55), .B1(n329), .B2(n354), .ZN(n80) );
  INV_X1 U73 ( .A(i[19]), .ZN(n354) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n368) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module register_file ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, 
        ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700,
         N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711,
         N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N1020,
         N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030,
         N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040,
         N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050,
         N1051, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3448, n3450,
         n3452, n3453, n3456, n3458, n3459, n3460, n3461, n3462, n3464, n3466,
         n3468, n3469, n3472, n3474, n3475, n3476, n3477, n3478, n3480, n3482,
         n3484, n3485, n3488, n3490, n3491, n3492, n3493, n3494, n3496, n3498,
         n3500, n3501, n3504, n3506, n3507, n3508, n3509, n3510, n3512, n3514,
         n3516, n3517, n3520, n3522, n3523, n3524, n3525, n3526, n3528, n3530,
         n3532, n3533, n3536, n3538, n3539, n3540, n3541, n3542, n3544, n3546,
         n3548, n3549, n3552, n3554, n3555, n3556, n3557, n3558, n3560, n3562,
         n3564, n3565, n3568, n3570, n3571, n3572, n3573, n3574, n3576, n3578,
         n3580, n3581, n3584, n3586, n3587, n3588, n3589, n3590, n3592, n3594,
         n3596, n3597, n3600, n3602, n3603, n3604, n3605, n3606, n3608, n3610,
         n3612, n3613, n3616, n3618, n3619, n3620, n3621, n3622, n3624, n3626,
         n3628, n3629, n3632, n3634, n3635, n3636, n3637, n3638, n3640, n3642,
         n3644, n3645, n3648, n3650, n3651, n3652, n3653, n3654, n3656, n3658,
         n3661, n3664, n3666, n3667, n3668, n3669, n3670, n3672, n3674, n3676,
         n3677, n3680, n3682, n3683, n3684, n3685, n3686, n3688, n3690, n3692,
         n3693, n3696, n3698, n3699, n3700, n3701, n3702, n3704, n3706, n3708,
         n3709, n3712, n3714, n3715, n3716, n3717, n3718, n3720, n3722, n3724,
         n3725, n3728, n3730, n3731, n3732, n3733, n3734, n3736, n3738, n3740,
         n3741, n3744, n3746, n3747, n3748, n3749, n3750, n3752, n3754, n3756,
         n3757, n3760, n3762, n3763, n3764, n3765, n3766, n3768, n3770, n3772,
         n3773, n3776, n3778, n3779, n3780, n3781, n3782, n3784, n3786, n3788,
         n3789, n3792, n3794, n3795, n3796, n3797, n3798, n3800, n3802, n3804,
         n3805, n3808, n3810, n3811, n3812, n3813, n3814, n3816, n3818, n3820,
         n3821, n3824, n3826, n3827, n3828, n3829, n3830, n3832, n3834, n3836,
         n3837, n3840, n3842, n3843, n3844, n3845, n3846, n3848, n3850, n3852,
         n3853, n3856, n3858, n3859, n3860, n3861, n3862, n3864, n3866, n3868,
         n3869, n3872, n3874, n3875, n3876, n3877, n3878, n3880, n3882, n3884,
         n3885, n3888, n3890, n3891, n3892, n3893, n3894, n3896, n3898, n3900,
         n3901, n3904, n3906, n3907, n3908, n3909, n3910, n3912, n3914, n3916,
         n3917, n3920, n3922, n3923, n3924, n3925, n3926, n3928, n3930, n3932,
         n3933, n3936, n3938, n3939, n3940, n3941, n3942, n3944, n3946, n3948,
         n3949, n3952, n3954, n3955, n3956, n3957, n3958, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n898, n899,
         n900, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n939, n940, n943, n954, n957, n959, n961,
         n970, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921;
  assign OUT1[0] = N690;
  assign OUT1[1] = N691;
  assign OUT1[2] = N692;
  assign OUT1[3] = N693;
  assign OUT1[4] = N694;
  assign OUT1[5] = N695;
  assign OUT1[6] = N696;
  assign OUT1[7] = N697;
  assign OUT1[8] = N698;
  assign OUT1[9] = N699;
  assign OUT1[10] = N700;
  assign OUT1[11] = N701;
  assign OUT1[12] = N702;
  assign OUT1[13] = N703;
  assign OUT1[14] = N704;
  assign OUT1[15] = N705;
  assign OUT1[16] = N706;
  assign OUT1[17] = N707;
  assign OUT1[18] = N708;
  assign OUT1[19] = N709;
  assign OUT1[20] = N710;
  assign OUT1[21] = N711;
  assign OUT1[22] = N712;
  assign OUT1[23] = N713;
  assign OUT1[24] = N714;
  assign OUT1[25] = N715;
  assign OUT1[26] = N716;
  assign OUT1[27] = N717;
  assign OUT1[28] = N718;
  assign OUT1[29] = N719;
  assign OUT1[30] = N720;
  assign OUT1[31] = N721;
  assign OUT2[0] = N1020;
  assign OUT2[1] = N1021;
  assign OUT2[2] = N1022;
  assign OUT2[3] = N1023;
  assign OUT2[4] = N1024;
  assign OUT2[5] = N1025;
  assign OUT2[6] = N1026;
  assign OUT2[7] = N1027;
  assign OUT2[8] = N1028;
  assign OUT2[9] = N1029;
  assign OUT2[10] = N1030;
  assign OUT2[11] = N1031;
  assign OUT2[12] = N1032;
  assign OUT2[13] = N1033;
  assign OUT2[14] = N1034;
  assign OUT2[15] = N1035;
  assign OUT2[16] = N1036;
  assign OUT2[17] = N1037;
  assign OUT2[18] = N1038;
  assign OUT2[19] = N1039;
  assign OUT2[20] = N1040;
  assign OUT2[21] = N1041;
  assign OUT2[22] = N1042;
  assign OUT2[23] = N1043;
  assign OUT2[24] = N1044;
  assign OUT2[25] = N1045;
  assign OUT2[26] = N1046;
  assign OUT2[27] = N1047;
  assign OUT2[28] = N1048;
  assign OUT2[29] = N1049;
  assign OUT2[30] = N1050;
  assign OUT2[31] = N1051;

  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n2901), .CK(CLK), .RN(n19056), .Q(
        n19905), .QN(n2364) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n2902), .CK(CLK), .RN(n19056), .Q(
        n19906), .QN(n2373) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n2903), .CK(CLK), .RN(n19056), .Q(
        n19907), .QN(n2382) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n2904), .CK(CLK), .RN(n19056), .Q(
        n19908), .QN(n2391) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n2905), .CK(CLK), .RN(n19056), .Q(
        n19909), .QN(n2400) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n2906), .CK(CLK), .RN(n19056), .Q(
        n19910), .QN(n2409) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n2907), .CK(CLK), .RN(n19056), .Q(n19911), .QN(n2418) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n2908), .CK(CLK), .RN(n19056), .Q(n19912), .QN(n2427) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n3069), .CK(CLK), .RN(n19056), .Q(
        n19255), .QN(n18210) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n3068), .CK(CLK), .RN(n19056), .Q(
        n19256), .QN(n18209) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n3067), .CK(CLK), .RN(n19056), .Q(
        n19257), .QN(n18208) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n3066), .CK(CLK), .RN(n19056), .Q(
        n19258), .QN(n18207) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n3065), .CK(CLK), .RN(n19056), .Q(
        n19259), .QN(n18206) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n3064), .CK(CLK), .RN(n19056), .Q(
        n19260), .QN(n18205) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n3063), .CK(CLK), .RN(n19056), .Q(
        n19261), .QN(n18204) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n3062), .CK(CLK), .RN(n19056), .Q(
        n19262), .QN(n18203) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n3005), .CK(CLK), .RN(n19056), .Q(
        n19215), .QN(n2218) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n3004), .CK(CLK), .RN(n19056), .Q(
        n19216), .QN(n2227) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n3003), .CK(CLK), .RN(n19056), .Q(
        n19217), .QN(n2236) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n3002), .CK(CLK), .RN(n19056), .Q(
        n19218), .QN(n2245) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n3001), .CK(CLK), .RN(n19056), .Q(
        n19219), .QN(n2254) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n3000), .CK(CLK), .RN(n19056), .Q(
        n19220), .QN(n2263) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n2999), .CK(CLK), .RN(n19056), .Q(
        n19221), .QN(n2272) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n2998), .CK(CLK), .RN(n19056), .Q(
        n19222), .QN(n2281) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n2973), .CK(CLK), .RN(n19056), .Q(
        n19239), .QN(n2219) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n2972), .CK(CLK), .RN(n19056), .Q(
        n19240), .QN(n2228) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n2971), .CK(CLK), .RN(n19056), .Q(
        n19241), .QN(n2237) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n2970), .CK(CLK), .RN(n19056), .Q(
        n19242), .QN(n2246) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n2969), .CK(CLK), .RN(n19056), .Q(
        n19243), .QN(n2255) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n2968), .CK(CLK), .RN(n19056), .Q(
        n19244), .QN(n2264) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n2967), .CK(CLK), .RN(n19056), .Q(
        n19245), .QN(n2273) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n2966), .CK(CLK), .RN(n19056), .Q(
        n19246), .QN(n2282) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n3813), .CK(CLK), .RN(n19056), .QN(
        n18076) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n9151), .CK(CLK), .RN(n19057), .Q(n19181), .QN(n2413) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n9055), .CK(CLK), .RN(n19056), .Q(n19285), .QN(n2421) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n3802), .CK(CLK), .RN(n19056), .Q(n19701), 
        .QN(n2419) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n3399), .CK(CLK), .RN(n19056), .QN(n18108) );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n2885), .CK(CLK), .RN(n19056), .Q(
        n19889), .QN(n2220) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n2886), .CK(CLK), .RN(n19056), .Q(
        n19890), .QN(n2229) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n2887), .CK(CLK), .RN(n19056), .Q(
        n19891), .QN(n2238) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n2888), .CK(CLK), .RN(n19056), .Q(
        n19892), .QN(n2247) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n2889), .CK(CLK), .RN(n19056), .Q(
        n19893), .QN(n2256) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n2890), .CK(CLK), .RN(n19056), .Q(
        n19894), .QN(n2265) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n2891), .CK(CLK), .RN(n19056), .Q(
        n19895), .QN(n2274) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n2892), .CK(CLK), .RN(n19056), .Q(
        n19896), .QN(n2283) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n2893), .CK(CLK), .RN(n19056), .Q(
        n19897), .QN(n2292) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n2894), .CK(CLK), .RN(n19056), .Q(
        n19898), .QN(n2301) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n2895), .CK(CLK), .RN(n19056), .Q(
        n19899), .QN(n2310) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n2896), .CK(CLK), .RN(n19056), .Q(
        n19900), .QN(n2319) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n2897), .CK(CLK), .RN(n19056), .Q(
        n19901), .QN(n2328) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n2898), .CK(CLK), .RN(n19056), .Q(
        n19902), .QN(n2337) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n2899), .CK(CLK), .RN(n19056), .Q(
        n19903), .QN(n2346) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n2900), .CK(CLK), .RN(n19056), .Q(
        n19904), .QN(n2355) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n2877), .CK(CLK), .RN(n19056), .Q(n19881), .QN(n2436) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n2878), .CK(CLK), .RN(n19056), .Q(n19882), .QN(n2445) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n2879), .CK(CLK), .RN(n19056), .Q(n19883), .QN(n2454) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n2880), .CK(CLK), .RN(n19056), .Q(n19884), .QN(n2463) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n2881), .CK(CLK), .RN(n19056), .Q(n19885), .QN(n2472) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n2882), .CK(CLK), .RN(n19056), .Q(n19886), .QN(n2481) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n2883), .CK(CLK), .RN(n19056), .Q(n19887), .QN(n2490) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n2884), .CK(CLK), .RN(n19056), .Q(n19888), .QN(n2499) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n3061), .CK(CLK), .RN(n19056), .Q(
        n19471), .QN(n17838) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n3060), .CK(CLK), .RN(n19056), .Q(
        n19472), .QN(n17837) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n3059), .CK(CLK), .RN(n19056), .Q(
        n19473), .QN(n17836) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n3058), .CK(CLK), .RN(n19056), .Q(
        n19474), .QN(n17835) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n3057), .CK(CLK), .RN(n19056), .Q(
        n19475), .QN(n17834) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n3055), .CK(CLK), .RN(n19056), .Q(
        n19477), .QN(n17832) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n3054), .CK(CLK), .RN(n19056), .Q(
        n19478), .QN(n17831) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n3053), .CK(CLK), .RN(n19056), .Q(
        n19479), .QN(n17830) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n3052), .CK(CLK), .RN(n19056), .Q(
        n19480), .QN(n17829) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n3051), .CK(CLK), .RN(n19056), .Q(
        n19481), .QN(n17828) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n3050), .CK(CLK), .RN(n19056), .Q(
        n19482), .QN(n17827) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n3049), .CK(CLK), .RN(n19056), .Q(
        n19483), .QN(n17826) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n3048), .CK(CLK), .RN(n19056), .Q(
        n19484), .QN(n17825) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n3047), .CK(CLK), .RN(n19056), .Q(n19485), .QN(n17824) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n3046), .CK(CLK), .RN(n19056), .Q(n19486), .QN(n17823) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n3045), .CK(CLK), .RN(n19056), .Q(n19487), .QN(n17822) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n3044), .CK(CLK), .RN(n19056), .Q(n19488), .QN(n17821) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n3043), .CK(CLK), .RN(n19056), .Q(n19489), .QN(n17820) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n3042), .CK(CLK), .RN(n19056), .Q(n19490), .QN(n17819) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n3041), .CK(CLK), .RN(n19056), .Q(n19491), .QN(n17818) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n3040), .CK(CLK), .RN(n19056), .Q(n19492), .QN(n17817) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n3039), .CK(CLK), .RN(n19056), .Q(n19493), .QN(n17816) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n3038), .CK(CLK), .RN(n19056), .Q(n19494), .QN(n17815) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n3175), .CK(CLK), .RN(n19056), .QN(
        n18180) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n3303), .CK(CLK), .RN(n19056), .QN(n18132) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n2997), .CK(CLK), .RN(n19056), .Q(
        n19343), .QN(n2290) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n2996), .CK(CLK), .RN(n19056), .Q(
        n19344), .QN(n2299) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n2995), .CK(CLK), .RN(n19056), .Q(
        n19345), .QN(n2308) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n2994), .CK(CLK), .RN(n19056), .Q(
        n19346), .QN(n2317) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n2993), .CK(CLK), .RN(n19056), .Q(
        n19347), .QN(n2326) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n2992), .CK(CLK), .RN(n19056), .Q(
        n19348), .QN(n2335) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n2991), .CK(CLK), .RN(n19056), .Q(
        n19349), .QN(n2344) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n2990), .CK(CLK), .RN(n19056), .Q(
        n19350), .QN(n2353) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n2989), .CK(CLK), .RN(n19056), .Q(
        n19351), .QN(n2362) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n2988), .CK(CLK), .RN(n19056), .Q(
        n19352), .QN(n2371) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n2987), .CK(CLK), .RN(n19056), .Q(
        n19353), .QN(n2380) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n2986), .CK(CLK), .RN(n19056), .Q(
        n19354), .QN(n2389) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n2985), .CK(CLK), .RN(n19056), .Q(
        n19355), .QN(n2398) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n2984), .CK(CLK), .RN(n19056), .Q(
        n19356), .QN(n2407) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n2983), .CK(CLK), .RN(n19056), .Q(n19357), .QN(n2416) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n2982), .CK(CLK), .RN(n19056), .Q(n19358), .QN(n2425) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n2981), .CK(CLK), .RN(n19056), .Q(n19359), .QN(n2434) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n2980), .CK(CLK), .RN(n19056), .Q(n19360), .QN(n2443) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n2979), .CK(CLK), .RN(n19056), .Q(n19361), .QN(n2452) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n2978), .CK(CLK), .RN(n19056), .Q(n19362), .QN(n2461) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n2977), .CK(CLK), .RN(n19056), .Q(n19363), .QN(n2470) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n2976), .CK(CLK), .RN(n19056), .Q(n19364), .QN(n2479) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n2975), .CK(CLK), .RN(n19056), .Q(n19365), .QN(n2488) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n2974), .CK(CLK), .RN(n19056), .Q(n19366), .QN(n2497) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n3808), .CK(CLK), .RN(n19056), .Q(n19797), .QN(n2414) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n18387), .CK(CLK), .RN(n19056), .Q(
        n19380), .QN(n2339) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n3804), .CK(CLK), .RN(n19056), .Q(n19389), 
        .QN(n2420) );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n3800), .CK(CLK), .RN(n19056), .Q(n19413), 
        .QN(n17943) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n2965), .CK(CLK), .RN(n19056), .Q(
        n19415), .QN(n2291) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n2964), .CK(CLK), .RN(n19056), .Q(
        n19416), .QN(n2300) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n2963), .CK(CLK), .RN(n19056), .Q(
        n19417), .QN(n2309) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n18386), .CK(CLK), .RN(n19056), .Q(
        n19418), .QN(n2318) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n2961), .CK(CLK), .RN(n19056), .Q(
        n19419), .QN(n2327) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n2960), .CK(CLK), .RN(n19056), .Q(
        n19420), .QN(n2336) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n2959), .CK(CLK), .RN(n19056), .Q(
        n19421), .QN(n2345) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n2958), .CK(CLK), .RN(n19056), .Q(
        n19422), .QN(n2354) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n2957), .CK(CLK), .RN(n19056), .Q(
        n19423), .QN(n2363) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n2956), .CK(CLK), .RN(n19056), .Q(
        n19424), .QN(n2372) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n2955), .CK(CLK), .RN(n19056), .Q(
        n19425), .QN(n2381) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n2954), .CK(CLK), .RN(n19056), .Q(
        n19426), .QN(n2390) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n2953), .CK(CLK), .RN(n19056), .Q(
        n19427), .QN(n2399) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n2952), .CK(CLK), .RN(n19056), .Q(
        n19428), .QN(n2408) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n2951), .CK(CLK), .RN(n19056), .Q(n19429), .QN(n2417) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n2950), .CK(CLK), .RN(n19056), .Q(n19430), .QN(n2426) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n2949), .CK(CLK), .RN(n19056), .Q(n19431), .QN(n2435) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n2948), .CK(CLK), .RN(n19056), .Q(n19432), .QN(n2444) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n2947), .CK(CLK), .RN(n19056), .Q(n19433), .QN(n2453) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n2946), .CK(CLK), .RN(n19056), .Q(n19434), .QN(n2462) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n2945), .CK(CLK), .RN(n19056), .Q(n19435), .QN(n2471) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n2944), .CK(CLK), .RN(n19056), .Q(n19436), .QN(n2480) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n2943), .CK(CLK), .RN(n19056), .Q(n19437), .QN(n2489) );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n2942), .CK(CLK), .RN(n19056), .Q(n19438), .QN(n2498) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n3079), .CK(CLK), .RN(n19056), .QN(
        n17904) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n3207), .CK(CLK), .RN(n19056), .QN(
        n17880) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n3335), .CK(CLK), .RN(n19056), .Q(n19453), 
        .QN(n17856) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n3143), .CK(CLK), .RN(n19056), .Q(n19509), .QN(n17800) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n3461), .CK(CLK), .RN(n19056), .QN(
        n18098) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n3829), .CK(CLK), .RN(n19056), .QN(
        n18075) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n3845), .CK(CLK), .RN(n19056), .QN(
        n18290) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n3861), .CK(CLK), .RN(n19056), .QN(
        n18289) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n3877), .CK(CLK), .RN(n19056), .QN(
        n18288) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n3893), .CK(CLK), .RN(n19056), .QN(
        n18287) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n3909), .CK(CLK), .RN(n19056), .QN(
        n18286) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n3456), .CK(CLK), .RN(n19056), .Q(
        n19775), .QN(n2216) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n3824), .CK(CLK), .RN(n19056), .Q(n19798), .QN(n2423) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n3840), .CK(CLK), .RN(n19056), .Q(n19639), .QN(n2432) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n3856), .CK(CLK), .RN(n19056), .Q(n19640), .QN(n2441) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n3872), .CK(CLK), .RN(n19056), .Q(n19641), .QN(n2450) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n3888), .CK(CLK), .RN(n19056), .Q(n19642), .QN(n2459) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n3904), .CK(CLK), .RN(n19056), .Q(n19643), .QN(n2468) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n9173), .CK(CLK), .RN(n19056), .Q(
        n19135), .QN(n2215) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n9150), .CK(CLK), .RN(n19057), .Q(n19182), .QN(n2422) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n9149), .CK(CLK), .RN(n19056), .Q(n19183), .QN(n2431) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n9148), .CK(CLK), .RN(n19056), .Q(n19184), .QN(n2440) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n9147), .CK(CLK), .RN(n19056), .Q(n19185), .QN(n2449) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n9146), .CK(CLK), .RN(n19056), .Q(n19186), .QN(n2458) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n9145), .CK(CLK), .RN(n19056), .Q(n19187), .QN(n2467) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n9077), .CK(CLK), .RN(n19056), .Q(
        n19191), .QN(n2223) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n9054), .CK(CLK), .RN(n19056), .Q(n19286), .QN(n2430) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n9053), .CK(CLK), .RN(n19056), .Q(n19287), .QN(n2439) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n9052), .CK(CLK), .RN(n19056), .Q(n19288), .QN(n2448) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n9051), .CK(CLK), .RN(n19056), .Q(n19289), .QN(n2457) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n9050), .CK(CLK), .RN(n19056), .Q(n19290), .QN(n2466) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n9049), .CK(CLK), .RN(n19056), .Q(n19291), .QN(n2475) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n3452), .CK(CLK), .RN(n19056), .Q(n19367), .QN(n2222) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n3820), .CK(CLK), .RN(n19056), .Q(n19390), 
        .QN(n2429) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n3836), .CK(CLK), .RN(n19056), .Q(n19223), 
        .QN(n2438) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n3852), .CK(CLK), .RN(n19056), .Q(n19224), 
        .QN(n2447) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n3868), .CK(CLK), .RN(n19056), .Q(n19225), 
        .QN(n2456) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n3884), .CK(CLK), .RN(n19056), .Q(n19226), 
        .QN(n2465) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n3900), .CK(CLK), .RN(n19056), .Q(n19227), 
        .QN(n2474) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n8986), .CK(CLK), .RN(n19056), .Q(n19338), 
        .QN(n18031) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n3101), .CK(CLK), .RN(n19056), .QN(
        n18234) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n3078), .CK(CLK), .RN(n19056), .QN(
        n17903) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n3077), .CK(CLK), .RN(n19056), .QN(
        n17902) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n3076), .CK(CLK), .RN(n19056), .QN(
        n17901) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n3075), .CK(CLK), .RN(n19056), .QN(
        n17900) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n3074), .CK(CLK), .RN(n19056), .QN(
        n17899) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n3073), .CK(CLK), .RN(n19056), .QN(
        n17898) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n3165), .CK(CLK), .RN(n19056), .Q(
        n19263), .QN(n18202) );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n3142), .CK(CLK), .RN(n19056), .Q(n19510), .QN(n17799) );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n3141), .CK(CLK), .RN(n19056), .Q(n19511), .QN(n17798) );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n3140), .CK(CLK), .RN(n19056), .Q(n19512), .QN(n17797) );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n3139), .CK(CLK), .RN(n19056), .Q(n19513), .QN(n17796) );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n3138), .CK(CLK), .RN(n19056), .Q(n19514), .QN(n17795) );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n3137), .CK(CLK), .RN(n19056), .Q(n19515), .QN(n17794) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n3197), .CK(CLK), .RN(n19056), .QN(
        n18322) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n3174), .CK(CLK), .RN(n19056), .QN(
        n18179) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n3173), .CK(CLK), .RN(n19056), .QN(
        n18178) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n3172), .CK(CLK), .RN(n19056), .QN(
        n18177) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n3171), .CK(CLK), .RN(n19056), .QN(
        n18176) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n3170), .CK(CLK), .RN(n19056), .QN(
        n18175) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n3169), .CK(CLK), .RN(n19056), .QN(
        n18174) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n3229), .CK(CLK), .RN(n19056), .QN(
        n18226) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n3206), .CK(CLK), .RN(n19056), .QN(
        n17879) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n3205), .CK(CLK), .RN(n19056), .QN(
        n17878) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n3204), .CK(CLK), .RN(n19056), .QN(
        n17877) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n3203), .CK(CLK), .RN(n19056), .QN(
        n17876) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n3202), .CK(CLK), .RN(n19056), .QN(
        n17875) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n3201), .CK(CLK), .RN(n19056), .QN(
        n17874) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n3325), .CK(CLK), .RN(n19056), .QN(
        n18306) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n3302), .CK(CLK), .RN(n19056), .QN(n18131) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n3301), .CK(CLK), .RN(n19056), .QN(n18130) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n3300), .CK(CLK), .RN(n19056), .QN(n18129) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n3299), .CK(CLK), .RN(n19056), .QN(n18128) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n3298), .CK(CLK), .RN(n19056), .QN(n18127) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n3297), .CK(CLK), .RN(n19056), .QN(n18126) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n3357), .CK(CLK), .RN(n19056), .Q(n19247), .QN(n18218) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n3334), .CK(CLK), .RN(n19056), .Q(n19454), 
        .QN(n17855) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n3333), .CK(CLK), .RN(n19056), .Q(n19455), 
        .QN(n17854) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n3332), .CK(CLK), .RN(n19056), .Q(n19456), 
        .QN(n17853) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n3331), .CK(CLK), .RN(n19056), .Q(n19457), 
        .QN(n17852) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n3330), .CK(CLK), .RN(n19056), .Q(n19458), 
        .QN(n17851) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n3329), .CK(CLK), .RN(n19056), .Q(n19459), 
        .QN(n17850) );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n3450), .CK(CLK), .RN(n19056), .Q(n19679), .QN(n2221) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n3818), .CK(CLK), .RN(n19056), .Q(n19702), 
        .QN(n2428) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n3834), .CK(CLK), .RN(n19056), .Q(n19607), 
        .QN(n2437) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n3850), .CK(CLK), .RN(n19056), .Q(n19608), 
        .QN(n2446) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n3866), .CK(CLK), .RN(n19056), .Q(n19609), 
        .QN(n2455) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n3882), .CK(CLK), .RN(n19056), .Q(n19610), 
        .QN(n2464) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n3898), .CK(CLK), .RN(n19056), .Q(n19611), 
        .QN(n2473) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n3421), .CK(CLK), .RN(n19056), .QN(
        n18298) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n3398), .CK(CLK), .RN(n19056), .QN(n18107) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n3397), .CK(CLK), .RN(n19056), .QN(n18106) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n3396), .CK(CLK), .RN(n19056), .QN(n18105) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n3395), .CK(CLK), .RN(n19056), .QN(n18104) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n3394), .CK(CLK), .RN(n19056), .QN(n18103) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n3393), .CK(CLK), .RN(n19056), .QN(n18102) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n3448), .CK(CLK), .RN(n19056), .Q(n19391), .QN(n17965) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n3816), .CK(CLK), .RN(n19056), .Q(n19414), 
        .QN(n17942) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n3832), .CK(CLK), .RN(n19056), .Q(n19231), 
        .QN(n18250) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n3848), .CK(CLK), .RN(n19056), .Q(n19232), 
        .QN(n18249) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n3864), .CK(CLK), .RN(n19056), .Q(n19233), 
        .QN(n18248) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n3880), .CK(CLK), .RN(n19056), .Q(n19234), 
        .QN(n18247) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n3896), .CK(CLK), .RN(n19056), .Q(n19235), 
        .QN(n18246) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n9205), .CK(CLK), .RN(n19056), .Q(
        n19463), .QN(n2217) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n3477), .CK(CLK), .RN(n19056), .QN(
        n18097) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n3493), .CK(CLK), .RN(n19056), .QN(
        n18096) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n3509), .CK(CLK), .RN(n19056), .QN(
        n18095) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n3525), .CK(CLK), .RN(n19056), .QN(
        n18094) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n3541), .CK(CLK), .RN(n19056), .QN(
        n18093) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n3557), .CK(CLK), .RN(n19056), .QN(
        n18092) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n3573), .CK(CLK), .RN(n19056), .QN(
        n18091) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n3589), .CK(CLK), .RN(n19056), .QN(
        n18090) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n3605), .CK(CLK), .RN(n19056), .QN(
        n18089) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n3621), .CK(CLK), .RN(n19056), .QN(
        n18088) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n3637), .CK(CLK), .RN(n19056), .QN(
        n18087) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n3653), .CK(CLK), .RN(n19056), .QN(
        n18086) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n3669), .CK(CLK), .RN(n19056), .QN(
        n18085) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n3685), .CK(CLK), .RN(n19056), .QN(
        n18084) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n3701), .CK(CLK), .RN(n19056), .QN(
        n18083) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n3717), .CK(CLK), .RN(n19056), .QN(
        n18082) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n3733), .CK(CLK), .RN(n19056), .QN(
        n18081) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n3749), .CK(CLK), .RN(n19056), .QN(
        n18080) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n3765), .CK(CLK), .RN(n19056), .QN(
        n18079) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n3781), .CK(CLK), .RN(n19056), .QN(
        n18078) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n3797), .CK(CLK), .RN(n19056), .QN(
        n18077) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n3925), .CK(CLK), .RN(n19056), .QN(
        n18285) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n3941), .CK(CLK), .RN(n19056), .QN(
        n18284) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n3957), .CK(CLK), .RN(n19056), .QN(
        n18283) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n3472), .CK(CLK), .RN(n19056), .Q(
        n19776), .QN(n2225) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n3488), .CK(CLK), .RN(n19056), .Q(
        n19777), .QN(n2234) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n3504), .CK(CLK), .RN(n19056), .Q(
        n19778), .QN(n2243) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n3520), .CK(CLK), .RN(n19056), .Q(
        n19779), .QN(n2252) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n3536), .CK(CLK), .RN(n19056), .Q(
        n19780), .QN(n2261) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n3552), .CK(CLK), .RN(n19056), .Q(
        n19781), .QN(n2270) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n3568), .CK(CLK), .RN(n19056), .Q(
        n19782), .QN(n2279) );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n3584), .CK(CLK), .RN(n19056), .Q(
        n19783), .QN(n2288) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n3600), .CK(CLK), .RN(n19056), .Q(
        n19784), .QN(n2297) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n3616), .CK(CLK), .RN(n19056), .Q(
        n19785), .QN(n2306) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n3632), .CK(CLK), .RN(n19056), .Q(
        n19786), .QN(n2315) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n3648), .CK(CLK), .RN(n19056), .Q(
        n19787), .QN(n2324) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n3664), .CK(CLK), .RN(n19056), .Q(
        n19788), .QN(n2333) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n3680), .CK(CLK), .RN(n19056), .Q(
        n19789), .QN(n2342) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n3696), .CK(CLK), .RN(n19056), .Q(
        n19790), .QN(n2351) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n3712), .CK(CLK), .RN(n19056), .Q(
        n19791), .QN(n2360) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n3728), .CK(CLK), .RN(n19056), .Q(
        n19792), .QN(n2369) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n3744), .CK(CLK), .RN(n19056), .Q(
        n19793), .QN(n2378) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n3760), .CK(CLK), .RN(n19056), .Q(
        n19794), .QN(n2387) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n3776), .CK(CLK), .RN(n19056), .Q(
        n19795), .QN(n2396) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n3792), .CK(CLK), .RN(n19056), .Q(
        n19796), .QN(n2405) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n3920), .CK(CLK), .RN(n19056), .Q(n19644), .QN(n2477) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n3936), .CK(CLK), .RN(n19056), .Q(n19645), .QN(n2486) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n3952), .CK(CLK), .RN(n19056), .Q(n19646), .QN(n2495) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n9172), .CK(CLK), .RN(n19056), .Q(
        n19136), .QN(n2224) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n9171), .CK(CLK), .RN(n19056), .Q(
        n19137), .QN(n2233) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n9170), .CK(CLK), .RN(n19056), .Q(
        n19138), .QN(n2242) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n9169), .CK(CLK), .RN(n19056), .Q(
        n19139), .QN(n2251) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n9168), .CK(CLK), .RN(n19056), .Q(
        n19140), .QN(n2260) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n9167), .CK(CLK), .RN(n19056), .Q(
        n19141), .QN(n2269) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n9166), .CK(CLK), .RN(n19056), .Q(
        n19142), .QN(n2278) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n9165), .CK(CLK), .RN(n19056), .Q(
        n19167), .QN(n2287) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n9164), .CK(CLK), .RN(n19056), .Q(
        n19168), .QN(n2296) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n9163), .CK(CLK), .RN(n19056), .Q(
        n19169), .QN(n2305) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n9162), .CK(CLK), .RN(n19056), .Q(
        n19170), .QN(n2314) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n9161), .CK(CLK), .RN(n19056), .Q(
        n19171), .QN(n2323) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n9160), .CK(CLK), .RN(n19056), .Q(
        n19172), .QN(n2332) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n9159), .CK(CLK), .RN(n19056), .Q(
        n19173), .QN(n2341) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n9158), .CK(CLK), .RN(n19056), .Q(
        n19174), .QN(n2350) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n9157), .CK(CLK), .RN(n19056), .Q(
        n19175), .QN(n2359) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n9156), .CK(CLK), .RN(n19056), .Q(
        n19176), .QN(n2368) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n9155), .CK(CLK), .RN(n19056), .Q(
        n19177), .QN(n2377) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n9154), .CK(CLK), .RN(n19056), .Q(
        n19178), .QN(n2386) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n9153), .CK(CLK), .RN(n19057), .Q(
        n19179), .QN(n2395) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n9152), .CK(CLK), .RN(n19057), .Q(
        n19180), .QN(n2404) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n9144), .CK(CLK), .RN(n19056), .Q(n19188), .QN(n2476) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n9143), .CK(CLK), .RN(n19056), .Q(n19189), .QN(n2485) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n9142), .CK(CLK), .RN(n19056), .Q(n19190), .QN(n2494) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n9076), .CK(CLK), .RN(n19056), .Q(
        n19192), .QN(n2232) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n9075), .CK(CLK), .RN(n19056), .Q(
        n19193), .QN(n2241) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n9074), .CK(CLK), .RN(n19056), .Q(
        n19194), .QN(n2250) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n9073), .CK(CLK), .RN(n19056), .Q(
        n19195), .QN(n2259) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n9072), .CK(CLK), .RN(n19056), .Q(
        n19196), .QN(n2268) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n9071), .CK(CLK), .RN(n19056), .Q(
        n19197), .QN(n2277) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n9070), .CK(CLK), .RN(n19056), .Q(
        n19198), .QN(n2286) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n9069), .CK(CLK), .RN(n19056), .Q(
        n19271), .QN(n2295) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n9068), .CK(CLK), .RN(n19056), .Q(
        n19272), .QN(n2304) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n9067), .CK(CLK), .RN(n19056), .Q(
        n19273), .QN(n2313) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n9066), .CK(CLK), .RN(n19056), .Q(
        n19274), .QN(n2322) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n9065), .CK(CLK), .RN(n19056), .Q(
        n19275), .QN(n2331) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n9064), .CK(CLK), .RN(n19056), .Q(
        n19276), .QN(n2340) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n9063), .CK(CLK), .RN(n19056), .Q(
        n19277), .QN(n2349) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n9062), .CK(CLK), .RN(n19056), .Q(
        n19278), .QN(n2358) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n9061), .CK(CLK), .RN(n19056), .Q(
        n19279), .QN(n2367) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n9060), .CK(CLK), .RN(n19056), .Q(
        n19280), .QN(n2376) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n9059), .CK(CLK), .RN(n19056), .Q(
        n19281), .QN(n2385) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n9058), .CK(CLK), .RN(n19056), .Q(
        n19282), .QN(n2394) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n9057), .CK(CLK), .RN(n19056), .Q(
        n19283), .QN(n2403) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n9056), .CK(CLK), .RN(n19056), .Q(
        n19284), .QN(n2412) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n9048), .CK(CLK), .RN(n19056), .Q(n19292), .QN(n2484) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n9047), .CK(CLK), .RN(n19056), .Q(n19293), .QN(n2493) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n9046), .CK(CLK), .RN(n19056), .Q(n19294), .QN(n2502) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n3629), .CK(CLK), .RN(n19056), .Q(
        n19306), .QN(n18063) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n3468), .CK(CLK), .RN(n19056), .Q(n19368), .QN(n2231) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n3484), .CK(CLK), .RN(n19056), .Q(n19369), .QN(n2240) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n3500), .CK(CLK), .RN(n19056), .Q(n19370), .QN(n2249) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n3516), .CK(CLK), .RN(n19056), .Q(n19371), .QN(n2258) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n3532), .CK(CLK), .RN(n19056), .Q(n19372), .QN(n2267) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n3548), .CK(CLK), .RN(n19056), .Q(n19373), .QN(n2276) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n3564), .CK(CLK), .RN(n19056), .Q(n19374), .QN(n2285) );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n3580), .CK(CLK), .RN(n19056), .Q(n19375), .QN(n2294) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n3596), .CK(CLK), .RN(n19056), .Q(n19376), .QN(n2303) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n3612), .CK(CLK), .RN(n19056), .Q(n19377), .QN(n2312) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n3628), .CK(CLK), .RN(n19056), .Q(n19378), .QN(n2321) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n3644), .CK(CLK), .RN(n19056), .Q(n19379), .QN(n2330) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n3676), .CK(CLK), .RN(n19056), .Q(n19381), .QN(n2348) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n3692), .CK(CLK), .RN(n19056), .Q(n19382), .QN(n2357) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n3708), .CK(CLK), .RN(n19056), .Q(n19383), .QN(n2366) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n3724), .CK(CLK), .RN(n19056), .Q(n19384), .QN(n2375) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n3740), .CK(CLK), .RN(n19056), .Q(n19385), .QN(n2384) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n3756), .CK(CLK), .RN(n19056), .Q(n19386), .QN(n2393) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n3772), .CK(CLK), .RN(n19056), .Q(n19387), .QN(n2402) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n3788), .CK(CLK), .RN(n19056), .Q(n19388), .QN(n2411) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n3916), .CK(CLK), .RN(n19056), .Q(n19228), 
        .QN(n2483) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n3932), .CK(CLK), .RN(n19056), .Q(n19229), 
        .QN(n2492) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n3948), .CK(CLK), .RN(n19056), .Q(n19230), 
        .QN(n2501) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n3658), .CK(CLK), .RN(n19056), .Q(n19692), .QN(n2338) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n9002), .CK(CLK), .RN(n19056), .Q(n19322), .QN(n18047) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n9000), .CK(CLK), .RN(n19056), .Q(n19324), .QN(n18045) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n8998), .CK(CLK), .RN(n19056), .Q(n19326), .QN(n18043) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n3056), .CK(CLK), .RN(n19056), .Q(
        n19476), .QN(n17833) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n3100), .CK(CLK), .RN(n19056), .QN(
        n18233) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n3099), .CK(CLK), .RN(n19056), .QN(
        n18232) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n3098), .CK(CLK), .RN(n19056), .QN(
        n18231) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n3097), .CK(CLK), .RN(n19056), .QN(
        n18230) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n3096), .CK(CLK), .RN(n19056), .QN(
        n18229) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n3095), .CK(CLK), .RN(n19056), .QN(
        n18228) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n3094), .CK(CLK), .RN(n19056), .QN(
        n18227) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n3093), .CK(CLK), .RN(n19056), .QN(
        n17918) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n3092), .CK(CLK), .RN(n19056), .QN(
        n17917) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n3091), .CK(CLK), .RN(n19056), .QN(
        n17916) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n3090), .CK(CLK), .RN(n19056), .QN(
        n17915) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n3089), .CK(CLK), .RN(n19056), .QN(
        n17914) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n3088), .CK(CLK), .RN(n19056), .QN(
        n17913) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n3087), .CK(CLK), .RN(n19056), .QN(
        n17912) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n3086), .CK(CLK), .RN(n19056), .QN(
        n17911) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n3085), .CK(CLK), .RN(n19056), .QN(
        n17910) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n3084), .CK(CLK), .RN(n19056), .QN(
        n17909) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n3083), .CK(CLK), .RN(n19056), .QN(
        n17908) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n3082), .CK(CLK), .RN(n19056), .QN(
        n17907) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n3081), .CK(CLK), .RN(n19056), .QN(
        n17906) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n3080), .CK(CLK), .RN(n19056), .QN(
        n17905) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n3072), .CK(CLK), .RN(n19056), .QN(
        n17897) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n3071), .CK(CLK), .RN(n19056), .QN(
        n17896) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n3070), .CK(CLK), .RN(n19056), .QN(
        n17895) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n3164), .CK(CLK), .RN(n19056), .Q(
        n19264), .QN(n18201) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n3163), .CK(CLK), .RN(n19056), .Q(
        n19265), .QN(n18200) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n3162), .CK(CLK), .RN(n19056), .Q(
        n19266), .QN(n18199) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n3161), .CK(CLK), .RN(n19056), .Q(
        n19267), .QN(n18198) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n3160), .CK(CLK), .RN(n19056), .Q(
        n19268), .QN(n18197) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n3159), .CK(CLK), .RN(n19056), .Q(
        n19269), .QN(n18196) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n3158), .CK(CLK), .RN(n19056), .Q(
        n19270), .QN(n18195) );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n3157), .CK(CLK), .RN(n19056), .Q(
        n19495), .QN(n17814) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n3156), .CK(CLK), .RN(n19056), .Q(
        n19496), .QN(n17813) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n3155), .CK(CLK), .RN(n19056), .Q(
        n19497), .QN(n17812) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n3154), .CK(CLK), .RN(n19056), .Q(
        n19498), .QN(n17811) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n3153), .CK(CLK), .RN(n19056), .Q(
        n19499), .QN(n17810) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n3152), .CK(CLK), .RN(n19056), .Q(
        n19500), .QN(n17809) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n3151), .CK(CLK), .RN(n19056), .Q(
        n19501), .QN(n17808) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n3150), .CK(CLK), .RN(n19056), .Q(
        n19502), .QN(n17807) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n3149), .CK(CLK), .RN(n19056), .Q(
        n19503), .QN(n17806) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n3148), .CK(CLK), .RN(n19056), .Q(
        n19504), .QN(n17805) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n3147), .CK(CLK), .RN(n19056), .Q(
        n19505), .QN(n17804) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n3146), .CK(CLK), .RN(n19056), .Q(
        n19506), .QN(n17803) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n3145), .CK(CLK), .RN(n19056), .Q(
        n19507), .QN(n17802) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n3144), .CK(CLK), .RN(n19056), .Q(
        n19508), .QN(n17801) );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n3136), .CK(CLK), .RN(n19056), .Q(n19516), .QN(n17793) );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n3135), .CK(CLK), .RN(n19056), .Q(n19517), .QN(n17792) );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n3134), .CK(CLK), .RN(n19056), .Q(n19518), .QN(n17791) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n3196), .CK(CLK), .RN(n19056), .QN(
        n18321) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n3195), .CK(CLK), .RN(n19056), .QN(
        n18320) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n3194), .CK(CLK), .RN(n19056), .QN(
        n18319) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n3193), .CK(CLK), .RN(n19056), .QN(
        n18318) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n3192), .CK(CLK), .RN(n19056), .QN(
        n18317) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n3191), .CK(CLK), .RN(n19056), .QN(
        n18316) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n3190), .CK(CLK), .RN(n19056), .QN(
        n18315) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n3189), .CK(CLK), .RN(n19056), .QN(
        n18194) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n3188), .CK(CLK), .RN(n19056), .QN(
        n18193) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n3187), .CK(CLK), .RN(n19056), .QN(
        n18192) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n3186), .CK(CLK), .RN(n19056), .QN(
        n18191) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n3185), .CK(CLK), .RN(n19056), .QN(
        n18190) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n3184), .CK(CLK), .RN(n19056), .QN(
        n18189) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n3183), .CK(CLK), .RN(n19056), .QN(
        n18188) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n3182), .CK(CLK), .RN(n19056), .QN(
        n18187) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n3181), .CK(CLK), .RN(n19056), .QN(
        n18186) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n3180), .CK(CLK), .RN(n19056), .QN(
        n18185) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n3179), .CK(CLK), .RN(n19056), .QN(
        n18184) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n3178), .CK(CLK), .RN(n19056), .QN(
        n18183) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n3177), .CK(CLK), .RN(n19056), .QN(
        n18182) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n3176), .CK(CLK), .RN(n19056), .QN(
        n18181) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n3168), .CK(CLK), .RN(n19056), .QN(
        n18173) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n3167), .CK(CLK), .RN(n19056), .QN(
        n18172) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n3166), .CK(CLK), .RN(n19056), .QN(
        n18171) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n3228), .CK(CLK), .RN(n19056), .QN(
        n18225) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n3227), .CK(CLK), .RN(n19056), .QN(
        n18224) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n3226), .CK(CLK), .RN(n19056), .QN(
        n18223) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n3225), .CK(CLK), .RN(n19056), .QN(
        n18222) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n3224), .CK(CLK), .RN(n19056), .QN(
        n18221) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n3223), .CK(CLK), .RN(n19056), .QN(
        n18220) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n3222), .CK(CLK), .RN(n19056), .QN(
        n18219) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n3221), .CK(CLK), .RN(n19056), .QN(
        n17894) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n3220), .CK(CLK), .RN(n19056), .QN(
        n17893) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n3219), .CK(CLK), .RN(n19056), .QN(
        n17892) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n3218), .CK(CLK), .RN(n19056), .QN(
        n17891) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n3217), .CK(CLK), .RN(n19056), .QN(
        n17890) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n3216), .CK(CLK), .RN(n19056), .QN(
        n17889) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n3215), .CK(CLK), .RN(n19056), .QN(
        n17888) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n3214), .CK(CLK), .RN(n19056), .QN(
        n17887) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n3213), .CK(CLK), .RN(n19056), .QN(
        n17886) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n3212), .CK(CLK), .RN(n19056), .QN(
        n17885) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n3211), .CK(CLK), .RN(n19056), .QN(
        n17884) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n3210), .CK(CLK), .RN(n19056), .QN(
        n17883) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n3209), .CK(CLK), .RN(n19056), .QN(
        n17882) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n3208), .CK(CLK), .RN(n19056), .QN(
        n17881) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n3200), .CK(CLK), .RN(n19056), .QN(
        n17873) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n3199), .CK(CLK), .RN(n19056), .QN(
        n17872) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n3198), .CK(CLK), .RN(n19056), .QN(
        n17871) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n3324), .CK(CLK), .RN(n19056), .QN(
        n18305) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n3323), .CK(CLK), .RN(n19056), .QN(
        n18304) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n3322), .CK(CLK), .RN(n19056), .QN(
        n18303) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n3321), .CK(CLK), .RN(n19056), .QN(
        n18302) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n3320), .CK(CLK), .RN(n19056), .QN(
        n18301) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n3319), .CK(CLK), .RN(n19056), .QN(
        n18300) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n3318), .CK(CLK), .RN(n19056), .QN(
        n18299) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n3317), .CK(CLK), .RN(n19056), .QN(
        n18146) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n3316), .CK(CLK), .RN(n19056), .QN(
        n18145) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n3315), .CK(CLK), .RN(n19056), .QN(
        n18144) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n3314), .CK(CLK), .RN(n19056), .QN(
        n18143) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n3313), .CK(CLK), .RN(n19056), .QN(
        n18142) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n3312), .CK(CLK), .RN(n19056), .QN(
        n18141) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n3311), .CK(CLK), .RN(n19056), .QN(
        n18140) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n3310), .CK(CLK), .RN(n19056), .QN(
        n18139) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n3309), .CK(CLK), .RN(n19056), .QN(
        n18138) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n3308), .CK(CLK), .RN(n19056), .QN(
        n18137) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n3307), .CK(CLK), .RN(n19056), .QN(
        n18136) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n3306), .CK(CLK), .RN(n19056), .QN(
        n18135) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n3305), .CK(CLK), .RN(n19056), .QN(
        n18134) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n3304), .CK(CLK), .RN(n19056), .QN(
        n18133) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n3296), .CK(CLK), .RN(n19056), .QN(n18125) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n3295), .CK(CLK), .RN(n19056), .QN(n18124) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n3294), .CK(CLK), .RN(n19056), .QN(n18123) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n3356), .CK(CLK), .RN(n19056), .Q(n19248), .QN(n18217) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n3355), .CK(CLK), .RN(n19056), .Q(n19249), .QN(n18216) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n3354), .CK(CLK), .RN(n19056), .Q(n19250), .QN(n18215) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n3353), .CK(CLK), .RN(n19056), .Q(n19251), .QN(n18214) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n3352), .CK(CLK), .RN(n19056), .Q(n19252), .QN(n18213) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n3351), .CK(CLK), .RN(n19056), .Q(n19253), .QN(n18212) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n3350), .CK(CLK), .RN(n19056), .Q(n19254), .QN(n18211) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n3349), .CK(CLK), .RN(n19056), .Q(n19439), .QN(n17870) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n3348), .CK(CLK), .RN(n19056), .Q(n19440), .QN(n17869) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n3347), .CK(CLK), .RN(n19056), .Q(n19441), .QN(n17868) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n3346), .CK(CLK), .RN(n19056), .Q(n19442), .QN(n17867) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n3345), .CK(CLK), .RN(n19056), .Q(n19443), .QN(n17866) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n3344), .CK(CLK), .RN(n19056), .Q(n19444), .QN(n17865) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n3343), .CK(CLK), .RN(n19056), .Q(n19445), .QN(n17864) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n3342), .CK(CLK), .RN(n19056), .Q(n19446), .QN(n17863) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n3341), .CK(CLK), .RN(n19056), .Q(n19447), .QN(n17862) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n3340), .CK(CLK), .RN(n19056), .Q(n19448), .QN(n17861) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n3339), .CK(CLK), .RN(n19056), .Q(n19449), .QN(n17860) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n3338), .CK(CLK), .RN(n19056), .Q(n19450), .QN(n17859) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n3337), .CK(CLK), .RN(n19056), .Q(n19451), .QN(n17858) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n3336), .CK(CLK), .RN(n19056), .Q(n19452), .QN(n17857) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n3328), .CK(CLK), .RN(n19056), .Q(n19460), 
        .QN(n17849) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n3327), .CK(CLK), .RN(n19056), .Q(n19461), 
        .QN(n17848) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n3326), .CK(CLK), .RN(n19056), .Q(n19462), 
        .QN(n17847) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n3466), .CK(CLK), .RN(n19056), .Q(n19680), .QN(n2230) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n3482), .CK(CLK), .RN(n19056), .Q(n19681), .QN(n2239) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n3498), .CK(CLK), .RN(n19056), .Q(n19682), .QN(n2248) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n3514), .CK(CLK), .RN(n19056), .Q(n19683), .QN(n2257) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n3530), .CK(CLK), .RN(n19056), .Q(n19684), .QN(n2266) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n3546), .CK(CLK), .RN(n19056), .Q(n19685), .QN(n2275) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n3562), .CK(CLK), .RN(n19056), .Q(n19686), .QN(n2284) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n3578), .CK(CLK), .RN(n19056), .Q(n19687), .QN(n2293) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n3594), .CK(CLK), .RN(n19056), .Q(n19688), .QN(n2302) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n3610), .CK(CLK), .RN(n19056), .Q(n19689), .QN(n2311) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n3626), .CK(CLK), .RN(n19056), .Q(n19690), .QN(n2320) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n3642), .CK(CLK), .RN(n19056), .Q(n19691), .QN(n2329) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n3674), .CK(CLK), .RN(n19056), .Q(n19693), .QN(n2347) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n3690), .CK(CLK), .RN(n19056), .Q(n19694), .QN(n2356) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n3706), .CK(CLK), .RN(n19056), .Q(n19695), .QN(n2365) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n3722), .CK(CLK), .RN(n19056), .Q(n19696), .QN(n2374) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n3738), .CK(CLK), .RN(n19056), .Q(n19697), .QN(n2383) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n3754), .CK(CLK), .RN(n19056), .Q(n19698), .QN(n2392) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n3770), .CK(CLK), .RN(n19056), .Q(n19699), .QN(n2401) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n3786), .CK(CLK), .RN(n19056), .Q(n19700), .QN(n2410) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n3914), .CK(CLK), .RN(n19056), .Q(n19612), 
        .QN(n2482) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n3930), .CK(CLK), .RN(n19056), .Q(n19613), 
        .QN(n2491) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n3946), .CK(CLK), .RN(n19056), .Q(n19614), 
        .QN(n2500) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n3381), .CK(CLK), .RN(n19056), .QN(
        n17979) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n3380), .CK(CLK), .RN(n19056), .QN(
        n17978) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n3379), .CK(CLK), .RN(n19056), .QN(
        n17977) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n3378), .CK(CLK), .RN(n19056), .QN(
        n17976) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n3377), .CK(CLK), .RN(n19056), .QN(
        n17975) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n3376), .CK(CLK), .RN(n19056), .QN(
        n17974) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n3375), .CK(CLK), .RN(n19056), .QN(
        n17973) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n3374), .CK(CLK), .RN(n19056), .QN(
        n17972) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n3373), .CK(CLK), .RN(n19056), .QN(
        n17971) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n3372), .CK(CLK), .RN(n19056), .QN(
        n17970) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n3371), .CK(CLK), .RN(n19056), .QN(
        n17969) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n3370), .CK(CLK), .RN(n19056), .QN(
        n17968) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n3369), .CK(CLK), .RN(n19056), .QN(
        n17967) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n3368), .CK(CLK), .RN(n19056), .QN(
        n17966) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n3420), .CK(CLK), .RN(n19056), .QN(
        n18297) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n3419), .CK(CLK), .RN(n19056), .QN(
        n18296) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n3418), .CK(CLK), .RN(n19056), .QN(
        n18295) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n3417), .CK(CLK), .RN(n19056), .QN(
        n18294) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n3416), .CK(CLK), .RN(n19056), .QN(
        n18293) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n3415), .CK(CLK), .RN(n19056), .QN(
        n18292) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n3414), .CK(CLK), .RN(n19056), .QN(
        n18291) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n3413), .CK(CLK), .RN(n19056), .QN(
        n18122) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n3412), .CK(CLK), .RN(n19056), .QN(
        n18121) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n3411), .CK(CLK), .RN(n19056), .QN(
        n18120) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n3410), .CK(CLK), .RN(n19056), .QN(
        n18119) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n3409), .CK(CLK), .RN(n19056), .QN(
        n18118) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n3408), .CK(CLK), .RN(n19056), .QN(
        n18117) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n3407), .CK(CLK), .RN(n19056), .QN(
        n18116) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n3406), .CK(CLK), .RN(n19056), .QN(
        n18115) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n3405), .CK(CLK), .RN(n19056), .QN(
        n18114) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n3404), .CK(CLK), .RN(n19056), .QN(
        n18113) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n3403), .CK(CLK), .RN(n19056), .QN(
        n18112) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n3402), .CK(CLK), .RN(n19056), .QN(
        n18111) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n3401), .CK(CLK), .RN(n19056), .QN(
        n18110) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n3400), .CK(CLK), .RN(n19056), .QN(
        n18109) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n3392), .CK(CLK), .RN(n19056), .QN(n18101) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n3391), .CK(CLK), .RN(n19056), .QN(n18100) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n3390), .CK(CLK), .RN(n19056), .QN(n18099) );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n3464), .CK(CLK), .RN(n19056), .Q(n19392), .QN(n17964) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n3480), .CK(CLK), .RN(n19056), .Q(n19393), .QN(n17963) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n3496), .CK(CLK), .RN(n19056), .Q(n19394), .QN(n17962) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n3512), .CK(CLK), .RN(n19056), .Q(n19395), .QN(n17961) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n3528), .CK(CLK), .RN(n19056), .Q(n19396), .QN(n17960) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n3544), .CK(CLK), .RN(n19056), .Q(n19397), .QN(n17959) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n3560), .CK(CLK), .RN(n19056), .Q(n19398), .QN(n17958) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n3576), .CK(CLK), .RN(n19056), .Q(n19399), .QN(n17957) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n3592), .CK(CLK), .RN(n19056), .Q(n19400), .QN(n17956) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n3608), .CK(CLK), .RN(n19056), .Q(n19401), .QN(n17955) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n3624), .CK(CLK), .RN(n19056), .Q(n19402), .QN(n17954) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n3640), .CK(CLK), .RN(n19056), .Q(n19403), .QN(n17953) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n3656), .CK(CLK), .RN(n19056), .Q(n19404), .QN(n17952) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n3672), .CK(CLK), .RN(n19056), .Q(n19405), .QN(n17951) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n3688), .CK(CLK), .RN(n19056), .Q(n19406), .QN(n17950) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n3704), .CK(CLK), .RN(n19056), .Q(n19407), .QN(n17949) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n3720), .CK(CLK), .RN(n19056), .Q(n19408), .QN(n17948) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n3736), .CK(CLK), .RN(n19056), .Q(n19409), .QN(n17947) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n3752), .CK(CLK), .RN(n19056), .Q(n19410), .QN(n17946) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n3768), .CK(CLK), .RN(n19056), .Q(n19411), .QN(n17945) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n3784), .CK(CLK), .RN(n19056), .Q(n19412), .QN(n17944) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n3912), .CK(CLK), .RN(n19056), .Q(n19236), 
        .QN(n18245) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n3928), .CK(CLK), .RN(n19056), .Q(n19237), 
        .QN(n18244) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n3944), .CK(CLK), .RN(n19056), .Q(n19238), 
        .QN(n18243) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n9183), .CK(CLK), .RN(n19056), .Q(n19533), .QN(n2415) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n9182), .CK(CLK), .RN(n19056), .Q(n19534), .QN(n2424) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n9181), .CK(CLK), .RN(n19056), .Q(n19535), .QN(n2433) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n9180), .CK(CLK), .RN(n19056), .Q(n19536), .QN(n2442) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n9179), .CK(CLK), .RN(n19056), .Q(n19537), .QN(n2451) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n9178), .CK(CLK), .RN(n19056), .Q(n19538), .QN(n2460) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n9177), .CK(CLK), .RN(n19056), .Q(n19539), .QN(n2469) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n9204), .CK(CLK), .RN(n19056), .Q(
        n19464), .QN(n2226) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n9203), .CK(CLK), .RN(n19056), .Q(
        n19465), .QN(n2235) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n9202), .CK(CLK), .RN(n19056), .Q(
        n19466), .QN(n2244) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n9201), .CK(CLK), .RN(n19056), .Q(
        n19467), .QN(n2253) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n9200), .CK(CLK), .RN(n19056), .Q(
        n19468), .QN(n2262) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n9199), .CK(CLK), .RN(n19056), .Q(
        n19469), .QN(n2271) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n9198), .CK(CLK), .RN(n19056), .Q(
        n19470), .QN(n2280) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n9197), .CK(CLK), .RN(n19056), .Q(
        n19519), .QN(n2289) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n9196), .CK(CLK), .RN(n19056), .Q(
        n19520), .QN(n2298) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n9195), .CK(CLK), .RN(n19056), .Q(
        n19521), .QN(n2307) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n9194), .CK(CLK), .RN(n19056), .Q(
        n19522), .QN(n2316) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n9193), .CK(CLK), .RN(n19056), .Q(
        n19523), .QN(n2325) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n9192), .CK(CLK), .RN(n19056), .Q(
        n19524), .QN(n2334) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n9191), .CK(CLK), .RN(n19056), .Q(
        n19525), .QN(n2343) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n9190), .CK(CLK), .RN(n19056), .Q(
        n19526), .QN(n2352) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n9189), .CK(CLK), .RN(n19056), .Q(
        n19527), .QN(n2361) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n9188), .CK(CLK), .RN(n19056), .Q(
        n19528), .QN(n2370) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n9187), .CK(CLK), .RN(n19056), .Q(
        n19529), .QN(n2379) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n9186), .CK(CLK), .RN(n19056), .Q(
        n19530), .QN(n2388) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n9185), .CK(CLK), .RN(n19056), .Q(
        n19531), .QN(n2397) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n9184), .CK(CLK), .RN(n19056), .Q(
        n19532), .QN(n2406) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n9176), .CK(CLK), .RN(n19056), .Q(n19540), .QN(n2478) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n9175), .CK(CLK), .RN(n19056), .Q(n19541), .QN(n2487) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n9174), .CK(CLK), .RN(n19056), .Q(n19542), .QN(n2496) );
  DFFR_X1 \REGISTERS_reg[0][7]  ( .D(n13849), .CK(CLK), .RN(n19056), .Q(n18385), .QN(n19127) );
  DFFR_X1 \REGISTERS_reg[0][6]  ( .D(n13850), .CK(CLK), .RN(n19056), .Q(n18384), .QN(n19128) );
  DFFR_X1 \REGISTERS_reg[0][5]  ( .D(n13851), .CK(CLK), .RN(n19056), .Q(n18383), .QN(n19129) );
  DFFR_X1 \REGISTERS_reg[0][4]  ( .D(n13852), .CK(CLK), .RN(n19056), .Q(n18382), .QN(n19130) );
  DFFR_X1 \REGISTERS_reg[0][3]  ( .D(n13853), .CK(CLK), .RN(n19056), .Q(n18381), .QN(n19131) );
  DFFR_X1 \REGISTERS_reg[0][2]  ( .D(n13854), .CK(CLK), .RN(n19056), .Q(n18380), .QN(n19132) );
  DFFR_X1 \REGISTERS_reg[0][1]  ( .D(n13855), .CK(CLK), .RN(n19056), .Q(n18379), .QN(n19133) );
  DFFR_X1 \REGISTERS_reg[0][0]  ( .D(n13856), .CK(CLK), .RN(n19056), .Q(n18378), .QN(n19134) );
  DFFR_X1 \REGISTERS_reg[0][31]  ( .D(n13825), .CK(CLK), .RN(n19056), .Q(
        n18369), .QN(n19143) );
  DFFR_X1 \REGISTERS_reg[0][30]  ( .D(n13826), .CK(CLK), .RN(n19056), .Q(
        n18368), .QN(n19144) );
  DFFR_X1 \REGISTERS_reg[0][29]  ( .D(n13827), .CK(CLK), .RN(n19056), .Q(
        n18367), .QN(n19145) );
  DFFR_X1 \REGISTERS_reg[0][28]  ( .D(n13828), .CK(CLK), .RN(n19056), .Q(
        n18366), .QN(n19146) );
  DFFR_X1 \REGISTERS_reg[0][27]  ( .D(n13829), .CK(CLK), .RN(n19056), .Q(
        n18365), .QN(n19147) );
  DFFR_X1 \REGISTERS_reg[0][26]  ( .D(n13830), .CK(CLK), .RN(n19056), .Q(
        n18364), .QN(n19148) );
  DFFR_X1 \REGISTERS_reg[0][25]  ( .D(n13831), .CK(CLK), .RN(n19056), .Q(
        n18363), .QN(n19149) );
  DFFR_X1 \REGISTERS_reg[0][24]  ( .D(n13832), .CK(CLK), .RN(n19056), .Q(
        n18362), .QN(n19150) );
  DFFR_X1 \REGISTERS_reg[0][23]  ( .D(n13833), .CK(CLK), .RN(n19056), .Q(
        n18361), .QN(n19151) );
  DFFR_X1 \REGISTERS_reg[0][22]  ( .D(n13834), .CK(CLK), .RN(n19056), .Q(
        n18360), .QN(n19152) );
  DFFR_X1 \REGISTERS_reg[0][21]  ( .D(n13835), .CK(CLK), .RN(n19056), .Q(
        n18359), .QN(n19153) );
  DFFR_X1 \REGISTERS_reg[0][20]  ( .D(n13836), .CK(CLK), .RN(n19056), .Q(
        n18358), .QN(n19154) );
  DFFR_X1 \REGISTERS_reg[0][19]  ( .D(n13837), .CK(CLK), .RN(n19056), .Q(
        n18357), .QN(n19155) );
  DFFR_X1 \REGISTERS_reg[0][18]  ( .D(n13838), .CK(CLK), .RN(n19056), .Q(
        n18356), .QN(n19156) );
  DFFR_X1 \REGISTERS_reg[0][17]  ( .D(n13839), .CK(CLK), .RN(n19056), .Q(
        n18355), .QN(n19157) );
  DFFR_X1 \REGISTERS_reg[0][16]  ( .D(n13840), .CK(CLK), .RN(n19056), .Q(
        n18354), .QN(n19158) );
  DFFR_X1 \REGISTERS_reg[0][15]  ( .D(n13841), .CK(CLK), .RN(n19056), .Q(
        n18353), .QN(n19159) );
  DFFR_X1 \REGISTERS_reg[0][14]  ( .D(n13842), .CK(CLK), .RN(n19056), .Q(
        n18352), .QN(n19160) );
  DFFR_X1 \REGISTERS_reg[0][13]  ( .D(n13843), .CK(CLK), .RN(n19056), .Q(
        n18351), .QN(n19161) );
  DFFR_X1 \REGISTERS_reg[0][12]  ( .D(n13844), .CK(CLK), .RN(n19056), .Q(
        n18350), .QN(n19162) );
  DFFR_X1 \REGISTERS_reg[0][11]  ( .D(n13845), .CK(CLK), .RN(n19056), .Q(
        n18349), .QN(n19163) );
  DFFR_X1 \REGISTERS_reg[0][10]  ( .D(n13846), .CK(CLK), .RN(n19056), .Q(
        n18348), .QN(n19164) );
  DFFR_X1 \REGISTERS_reg[0][9]  ( .D(n13847), .CK(CLK), .RN(n19056), .Q(n18347), .QN(n19165) );
  DFFR_X1 \REGISTERS_reg[0][8]  ( .D(n13848), .CK(CLK), .RN(n19056), .Q(n18346), .QN(n19166) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n3811), .CK(CLK), .RN(n19056), .Q(n17728), .QN(n19581) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n3805), .CK(CLK), .RN(n19056), .Q(n18052), .QN(n19317) );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n9023), .CK(CLK), .RN(n19056), .Q(n17712), 
        .QN(n19597) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n8991), .CK(CLK), .RN(n19056), .Q(n18036), 
        .QN(n19333) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n3271), .CK(CLK), .RN(n19056), .Q(n17584), .QN(n19717) );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n3812), .CK(CLK), .RN(n19056), .QN(
        n19749) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n3111), .CK(CLK), .RN(n19056), .QN(
        n19765) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n3239), .CK(CLK), .RN(n19056), .Q(n17536), .QN(n19813) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n3367), .CK(CLK), .RN(n19056), .QN(n19823) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n3814), .CK(CLK), .RN(n19056), .Q(n17504), .QN(n19855) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n3810), .CK(CLK), .RN(n19056), .Q(n17480), .QN(n19879) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n3462), .CK(CLK), .RN(n19056), .Q(
        n17526), .QN(n19833) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n3830), .CK(CLK), .RN(n19056), .Q(n17503), .QN(n19856) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n3846), .CK(CLK), .RN(n19056), .Q(n17662), .QN(n19663) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n3862), .CK(CLK), .RN(n19056), .Q(n17661), .QN(n19664) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n3878), .CK(CLK), .RN(n19056), .Q(n17660), .QN(n19665) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n3894), .CK(CLK), .RN(n19056), .Q(n17659), .QN(n19666) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n3910), .CK(CLK), .RN(n19056), .Q(n17658), .QN(n19667) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n3460), .CK(CLK), .RN(n19056), .QN(
        n19727) );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n3828), .CK(CLK), .RN(n19056), .QN(
        n19750) );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n3844), .CK(CLK), .RN(n19056), .QN(
        n19623) );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n3860), .CK(CLK), .RN(n19056), .QN(
        n19624) );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n3876), .CK(CLK), .RN(n19056), .QN(
        n19625) );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n3892), .CK(CLK), .RN(n19056), .QN(
        n19626) );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n3908), .CK(CLK), .RN(n19056), .QN(
        n19627) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n3459), .CK(CLK), .RN(n19056), .Q(
        n17750), .QN(n19559) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n3827), .CK(CLK), .RN(n19056), .Q(n17727), .QN(n19582) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n3843), .CK(CLK), .RN(n19056), .Q(n17766), .QN(n19543) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n3859), .CK(CLK), .RN(n19056), .Q(n17765), .QN(n19544) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n3875), .CK(CLK), .RN(n19056), .Q(n17764), .QN(n19545) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n3891), .CK(CLK), .RN(n19056), .Q(n17763), .QN(n19546) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n3907), .CK(CLK), .RN(n19056), .Q(n17762), .QN(n19547) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n3458), .CK(CLK), .RN(n19056), .Q(
        n17502), .QN(n19857) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n3826), .CK(CLK), .RN(n19056), .Q(n17479), .QN(n19880) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n3842), .CK(CLK), .RN(n19056), .Q(n17654), .QN(n19671) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n3858), .CK(CLK), .RN(n19056), .Q(n17653), .QN(n19672) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n3874), .CK(CLK), .RN(n19056), .Q(n17652), .QN(n19673) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n3890), .CK(CLK), .RN(n19056), .Q(n17651), .QN(n19674) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n3906), .CK(CLK), .RN(n19056), .Q(n17650), .QN(n19675) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n3453), .CK(CLK), .RN(n19056), .Q(
        n18074), .QN(n19295) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n3821), .CK(CLK), .RN(n19056), .Q(n18051), .QN(n19318) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n3837), .CK(CLK), .RN(n19056), .Q(n18282), .QN(n19199) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n3853), .CK(CLK), .RN(n19056), .Q(n18281), .QN(n19200) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n3869), .CK(CLK), .RN(n19056), .Q(n18280), .QN(n19201) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n3885), .CK(CLK), .RN(n19056), .Q(n18279), .QN(n19202) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n3901), .CK(CLK), .RN(n19056), .Q(n18278), .QN(n19203) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n9045), .CK(CLK), .RN(n19056), .Q(n17758), .QN(n19551) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n9022), .CK(CLK), .RN(n19056), .Q(n17711), 
        .QN(n19598) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n9021), .CK(CLK), .RN(n19056), .Q(n17710), 
        .QN(n19599) );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n9020), .CK(CLK), .RN(n19056), .Q(n17709), 
        .QN(n19600) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n9019), .CK(CLK), .RN(n19056), .Q(n17708), 
        .QN(n19601) );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n9018), .CK(CLK), .RN(n19056), .Q(n17707), 
        .QN(n19602) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n9017), .CK(CLK), .RN(n19056), .Q(n17706), 
        .QN(n19603) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n9013), .CK(CLK), .RN(n19056), .Q(n18274), .QN(n19207) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n8990), .CK(CLK), .RN(n19056), .Q(n18035), 
        .QN(n19334) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n8989), .CK(CLK), .RN(n19056), .Q(n18034), 
        .QN(n19335) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n8988), .CK(CLK), .RN(n19056), .Q(n18033), 
        .QN(n19336) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n8987), .CK(CLK), .RN(n19056), .Q(n18032), 
        .QN(n19337) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n8985), .CK(CLK), .RN(n19056), .Q(n18030), 
        .QN(n19339) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n3133), .CK(CLK), .RN(n19056), .QN(
        n19631) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n3110), .CK(CLK), .RN(n19056), .QN(
        n19766) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n3109), .CK(CLK), .RN(n19056), .QN(
        n19767) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n3108), .CK(CLK), .RN(n19056), .QN(
        n19768) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n3107), .CK(CLK), .RN(n19056), .QN(
        n19769) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n3106), .CK(CLK), .RN(n19056), .QN(
        n19770) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n3105), .CK(CLK), .RN(n19056), .QN(
        n19771) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n3261), .CK(CLK), .RN(n19056), .Q(
        n17670), .QN(n19647) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n3238), .CK(CLK), .RN(n19056), .Q(n17535), .QN(n19814) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n3237), .CK(CLK), .RN(n19056), .Q(n17534), .QN(n19815) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n3236), .CK(CLK), .RN(n19056), .Q(n17533), .QN(n19816) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n3235), .CK(CLK), .RN(n19056), .Q(n17532), .QN(n19817) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n3234), .CK(CLK), .RN(n19056), .Q(n17531), .QN(n19818) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n3233), .CK(CLK), .RN(n19056), .Q(n17530), .QN(n19819) );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n3293), .CK(CLK), .RN(n19056), .Q(
        n17686), .QN(n19615) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n3270), .CK(CLK), .RN(n19056), .Q(n17583), .QN(n19718) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n3269), .CK(CLK), .RN(n19056), .Q(n17582), .QN(n19719) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n3268), .CK(CLK), .RN(n19056), .Q(n17581), .QN(n19720) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n3267), .CK(CLK), .RN(n19056), .Q(n17580), .QN(n19721) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n3266), .CK(CLK), .RN(n19056), .Q(n17579), .QN(n19722) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n3265), .CK(CLK), .RN(n19056), .Q(n17578), .QN(n19723) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n3389), .CK(CLK), .RN(n19056), .QN(
        n19655) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n3366), .CK(CLK), .RN(n19056), .QN(n19824) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n3365), .CK(CLK), .RN(n19056), .QN(n19825) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n3364), .CK(CLK), .RN(n19056), .QN(n19826) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n3363), .CK(CLK), .RN(n19056), .QN(n19827) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n3362), .CK(CLK), .RN(n19056), .QN(n19828) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n3361), .CK(CLK), .RN(n19056), .QN(n19829) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n19107), .CK(CLK), .RN(n19056), .Q(
        n17694) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n19109), .CK(CLK), .RN(n19056), .Q(
        n17693) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n19111), .CK(CLK), .RN(n19056), .Q(
        n17692) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n19113), .CK(CLK), .RN(n19056), .Q(
        n17691) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n19115), .CK(CLK), .RN(n19056), .Q(
        n17690) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n19117), .CK(CLK), .RN(n19056), .Q(
        n17689) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n19119), .CK(CLK), .RN(n19056), .Q(
        n17688) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n19121), .CK(CLK), .RN(n19056), .Q(
        n17687) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n3478), .CK(CLK), .RN(n19056), .Q(
        n17525), .QN(n19834) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n3494), .CK(CLK), .RN(n19056), .Q(
        n17524), .QN(n19835) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n3510), .CK(CLK), .RN(n19056), .Q(
        n17523), .QN(n19836) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n3526), .CK(CLK), .RN(n19056), .Q(
        n17522), .QN(n19837) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n3542), .CK(CLK), .RN(n19056), .Q(
        n17521), .QN(n19838) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n3558), .CK(CLK), .RN(n19056), .Q(
        n17520), .QN(n19839) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n3574), .CK(CLK), .RN(n19056), .Q(
        n17519), .QN(n19840) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n3590), .CK(CLK), .RN(n19056), .Q(
        n17518), .QN(n19841) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n3606), .CK(CLK), .RN(n19056), .Q(
        n17517), .QN(n19842) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n3622), .CK(CLK), .RN(n19056), .Q(
        n17516), .QN(n19843) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n3638), .CK(CLK), .RN(n19056), .Q(
        n17515), .QN(n19844) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n3654), .CK(CLK), .RN(n19056), .Q(
        n17514), .QN(n19845) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n3670), .CK(CLK), .RN(n19056), .Q(
        n17513), .QN(n19846) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n3686), .CK(CLK), .RN(n19056), .Q(
        n17512), .QN(n19847) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n3702), .CK(CLK), .RN(n19056), .Q(
        n17511), .QN(n19848) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n3718), .CK(CLK), .RN(n19056), .Q(
        n17510), .QN(n19849) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n3734), .CK(CLK), .RN(n19056), .Q(
        n17509), .QN(n19850) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n3750), .CK(CLK), .RN(n19056), .Q(
        n17508), .QN(n19851) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n3766), .CK(CLK), .RN(n19056), .Q(
        n17507), .QN(n19852) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n3782), .CK(CLK), .RN(n19056), .Q(
        n17506), .QN(n19853) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n3798), .CK(CLK), .RN(n19056), .Q(
        n17505), .QN(n19854) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n3926), .CK(CLK), .RN(n19056), .Q(n17657), .QN(n19668) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n3942), .CK(CLK), .RN(n19056), .Q(n17656), .QN(n19669) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n3958), .CK(CLK), .RN(n19056), .Q(n17655), .QN(n19670) );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n3476), .CK(CLK), .RN(n19056), .QN(
        n19728) );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n3492), .CK(CLK), .RN(n19056), .QN(
        n19729) );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n3508), .CK(CLK), .RN(n19056), .QN(
        n19730) );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n3524), .CK(CLK), .RN(n19056), .QN(
        n19731) );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n3540), .CK(CLK), .RN(n19056), .QN(
        n19732) );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n3556), .CK(CLK), .RN(n19056), .QN(
        n19733) );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n3572), .CK(CLK), .RN(n19056), .QN(
        n19734) );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n3588), .CK(CLK), .RN(n19056), .QN(
        n19735) );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n3604), .CK(CLK), .RN(n19056), .QN(
        n19736) );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n3620), .CK(CLK), .RN(n19056), .QN(
        n19737) );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n3636), .CK(CLK), .RN(n19056), .QN(
        n19738) );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n3652), .CK(CLK), .RN(n19056), .QN(
        n19739) );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n3668), .CK(CLK), .RN(n19056), .QN(
        n19740) );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n3684), .CK(CLK), .RN(n19056), .QN(
        n19741) );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n3700), .CK(CLK), .RN(n19056), .QN(
        n19742) );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n3716), .CK(CLK), .RN(n19056), .QN(
        n19743) );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n3732), .CK(CLK), .RN(n19056), .QN(
        n19744) );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n3748), .CK(CLK), .RN(n19056), .QN(
        n19745) );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n3764), .CK(CLK), .RN(n19056), .QN(
        n19746) );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n3780), .CK(CLK), .RN(n19056), .QN(
        n19747) );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n3796), .CK(CLK), .RN(n19056), .QN(
        n19748) );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n3924), .CK(CLK), .RN(n19056), .QN(
        n19628) );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n3940), .CK(CLK), .RN(n19056), .QN(
        n19629) );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n3956), .CK(CLK), .RN(n19056), .QN(
        n19630) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n3475), .CK(CLK), .RN(n19056), .Q(
        n17749), .QN(n19560) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n3491), .CK(CLK), .RN(n19056), .Q(
        n17748), .QN(n19561) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n3507), .CK(CLK), .RN(n19056), .Q(
        n17747), .QN(n19562) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n3523), .CK(CLK), .RN(n19056), .Q(
        n17746), .QN(n19563) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n3539), .CK(CLK), .RN(n19056), .Q(
        n17745), .QN(n19564) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n3555), .CK(CLK), .RN(n19056), .Q(
        n17744), .QN(n19565) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n3571), .CK(CLK), .RN(n19056), .Q(
        n17743), .QN(n19566) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n3587), .CK(CLK), .RN(n19056), .Q(
        n17742), .QN(n19567) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n3603), .CK(CLK), .RN(n19056), .Q(
        n17741), .QN(n19568) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n3619), .CK(CLK), .RN(n19056), .Q(
        n17740), .QN(n19569) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n3635), .CK(CLK), .RN(n19056), .Q(
        n17739), .QN(n19570) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n3651), .CK(CLK), .RN(n19056), .Q(
        n17738), .QN(n19571) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n3667), .CK(CLK), .RN(n19056), .Q(
        n17737), .QN(n19572) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n3683), .CK(CLK), .RN(n19056), .Q(
        n17736), .QN(n19573) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n3699), .CK(CLK), .RN(n19056), .Q(
        n17735), .QN(n19574) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n3715), .CK(CLK), .RN(n19056), .Q(
        n17734), .QN(n19575) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n3731), .CK(CLK), .RN(n19056), .Q(
        n17733), .QN(n19576) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n3747), .CK(CLK), .RN(n19056), .Q(
        n17732), .QN(n19577) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n3763), .CK(CLK), .RN(n19056), .Q(
        n17731), .QN(n19578) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n3779), .CK(CLK), .RN(n19056), .Q(
        n17730), .QN(n19579) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n3795), .CK(CLK), .RN(n19056), .Q(
        n17729), .QN(n19580) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n3923), .CK(CLK), .RN(n19056), .Q(n17761), .QN(n19548) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n3939), .CK(CLK), .RN(n19056), .Q(n17760), .QN(n19549) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n3955), .CK(CLK), .RN(n19056), .Q(n17759), .QN(n19550) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n3474), .CK(CLK), .RN(n19056), .Q(
        n17501), .QN(n19858) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n3490), .CK(CLK), .RN(n19056), .Q(
        n17500), .QN(n19859) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n3506), .CK(CLK), .RN(n19056), .Q(
        n17499), .QN(n19860) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n3522), .CK(CLK), .RN(n19056), .Q(
        n17498), .QN(n19861) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n3538), .CK(CLK), .RN(n19056), .Q(
        n17497), .QN(n19862) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n3554), .CK(CLK), .RN(n19056), .Q(
        n17496), .QN(n19863) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n3570), .CK(CLK), .RN(n19056), .Q(
        n17495), .QN(n19864) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n3586), .CK(CLK), .RN(n19056), .Q(
        n17494), .QN(n19865) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n3602), .CK(CLK), .RN(n19056), .Q(
        n17493), .QN(n19866) );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n3618), .CK(CLK), .RN(n19056), .Q(
        n17492), .QN(n19867) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n3634), .CK(CLK), .RN(n19056), .Q(
        n17491), .QN(n19868) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n3650), .CK(CLK), .RN(n19056), .Q(
        n17490), .QN(n19869) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n3666), .CK(CLK), .RN(n19056), .Q(
        n17489), .QN(n19870) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n3682), .CK(CLK), .RN(n19056), .Q(
        n17488), .QN(n19871) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n3698), .CK(CLK), .RN(n19056), .Q(
        n17487), .QN(n19872) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n3714), .CK(CLK), .RN(n19056), .Q(
        n17486), .QN(n19873) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n3730), .CK(CLK), .RN(n19056), .Q(
        n17485), .QN(n19874) );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n3746), .CK(CLK), .RN(n19056), .Q(
        n17484), .QN(n19875) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n3762), .CK(CLK), .RN(n19056), .Q(
        n17483), .QN(n19876) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n3778), .CK(CLK), .RN(n19056), .Q(
        n17482), .QN(n19877) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n3794), .CK(CLK), .RN(n19056), .Q(
        n17481), .QN(n19878) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n3922), .CK(CLK), .RN(n19056), .Q(n17649), .QN(n19676) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n3938), .CK(CLK), .RN(n19056), .Q(n17648), .QN(n19677) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n3954), .CK(CLK), .RN(n19056), .Q(n17647), .QN(n19678) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n3469), .CK(CLK), .RN(n19056), .Q(
        n18073), .QN(n19296) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n3485), .CK(CLK), .RN(n19056), .Q(
        n18072), .QN(n19297) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n3501), .CK(CLK), .RN(n19056), .Q(
        n18071), .QN(n19298) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n3517), .CK(CLK), .RN(n19056), .Q(
        n18070), .QN(n19299) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n3533), .CK(CLK), .RN(n19056), .Q(
        n18069), .QN(n19300) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n3549), .CK(CLK), .RN(n19056), .Q(
        n18068), .QN(n19301) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n3565), .CK(CLK), .RN(n19056), .Q(
        n18067), .QN(n19302) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n3581), .CK(CLK), .RN(n19056), .Q(
        n18066), .QN(n19303) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n3597), .CK(CLK), .RN(n19056), .Q(
        n18065), .QN(n19304) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n3613), .CK(CLK), .RN(n19056), .Q(
        n18064), .QN(n19305) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n3645), .CK(CLK), .RN(n19056), .Q(
        n18062), .QN(n19307) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n3661), .CK(CLK), .RN(n19056), .Q(
        n18061), .QN(n19308) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n3677), .CK(CLK), .RN(n19056), .Q(
        n18060), .QN(n19309) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n3693), .CK(CLK), .RN(n19056), .Q(
        n18059), .QN(n19310) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n3709), .CK(CLK), .RN(n19056), .Q(
        n18058), .QN(n19311) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n3725), .CK(CLK), .RN(n19056), .Q(
        n18057), .QN(n19312) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n3741), .CK(CLK), .RN(n19056), .Q(
        n18056), .QN(n19313) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n3757), .CK(CLK), .RN(n19056), .Q(
        n18055), .QN(n19314) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n3773), .CK(CLK), .RN(n19056), .Q(
        n18054), .QN(n19315) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n3789), .CK(CLK), .RN(n19056), .Q(
        n18053), .QN(n19316) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n3917), .CK(CLK), .RN(n19056), .Q(n18277), .QN(n19204) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n3933), .CK(CLK), .RN(n19056), .Q(n18276), .QN(n19205) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n3949), .CK(CLK), .RN(n19056), .Q(n18275), .QN(n19206) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n9044), .CK(CLK), .RN(n19056), .Q(n17757), .QN(n19552) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n9043), .CK(CLK), .RN(n19056), .Q(n17756), .QN(n19553) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n9042), .CK(CLK), .RN(n19056), .Q(n17755), .QN(n19554) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n9041), .CK(CLK), .RN(n19056), .Q(n17754), .QN(n19555) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n9040), .CK(CLK), .RN(n19056), .Q(n17753), .QN(n19556) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n9039), .CK(CLK), .RN(n19056), .Q(n17752), .QN(n19557) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n9038), .CK(CLK), .RN(n19056), .Q(n17751), .QN(n19558) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n9037), .CK(CLK), .RN(n19056), .Q(n17726), .QN(n19583) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n9036), .CK(CLK), .RN(n19056), .Q(n17725), .QN(n19584) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n9035), .CK(CLK), .RN(n19056), .Q(n17724), .QN(n19585) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n9034), .CK(CLK), .RN(n19056), .Q(n17723), .QN(n19586) );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n9033), .CK(CLK), .RN(n19056), .Q(n17722), .QN(n19587) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n9032), .CK(CLK), .RN(n19056), .Q(n17721), .QN(n19588) );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n9031), .CK(CLK), .RN(n19056), .Q(n17720), .QN(n19589) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n9030), .CK(CLK), .RN(n19056), .Q(n17719), .QN(n19590) );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n9029), .CK(CLK), .RN(n19056), .Q(n17718), .QN(n19591) );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n9028), .CK(CLK), .RN(n19056), .Q(n17717), .QN(n19592) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n9027), .CK(CLK), .RN(n19056), .Q(n17716), .QN(n19593) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n9026), .CK(CLK), .RN(n19056), .Q(n17715), .QN(n19594) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n9025), .CK(CLK), .RN(n19056), .Q(n17714), .QN(n19595) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n9024), .CK(CLK), .RN(n19056), .Q(n17713), .QN(n19596) );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n9016), .CK(CLK), .RN(n19056), .Q(n17705), 
        .QN(n19604) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n9015), .CK(CLK), .RN(n19056), .Q(n17704), 
        .QN(n19605) );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n9014), .CK(CLK), .RN(n19056), .Q(n17703), 
        .QN(n19606) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n9012), .CK(CLK), .RN(n19056), .Q(n18273), .QN(n19208) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n9011), .CK(CLK), .RN(n19056), .Q(n18272), .QN(n19209) );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n9010), .CK(CLK), .RN(n19056), .Q(n18271), .QN(n19210) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n9009), .CK(CLK), .RN(n19056), .Q(n18270), .QN(n19211) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n9008), .CK(CLK), .RN(n19056), .Q(n18269), .QN(n19212) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n9007), .CK(CLK), .RN(n19056), .Q(n18268), .QN(n19213) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n9006), .CK(CLK), .RN(n19056), .Q(n18267), .QN(n19214) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n9005), .CK(CLK), .RN(n19056), .Q(n18050), .QN(n19319) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n9004), .CK(CLK), .RN(n19056), .Q(n18049), .QN(n19320) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n9003), .CK(CLK), .RN(n19056), .Q(n18048), .QN(n19321) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n9001), .CK(CLK), .RN(n19056), .Q(n18046), .QN(n19323) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n8999), .CK(CLK), .RN(n19056), .Q(n18044), .QN(n19325) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n8997), .CK(CLK), .RN(n19056), .Q(n18042), .QN(n19327) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n8996), .CK(CLK), .RN(n19056), .Q(n18041), .QN(n19328) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n8995), .CK(CLK), .RN(n19056), .Q(n18040), .QN(n19329) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n8994), .CK(CLK), .RN(n19056), .Q(n18039), .QN(n19330) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n8993), .CK(CLK), .RN(n19056), .Q(n18038), .QN(n19331) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n8992), .CK(CLK), .RN(n19056), .Q(n18037), .QN(n19332) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n8984), .CK(CLK), .RN(n19056), .Q(n18029), 
        .QN(n19340) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n8983), .CK(CLK), .RN(n19056), .Q(n18028), 
        .QN(n19341) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n8982), .CK(CLK), .RN(n19056), .Q(n18027), 
        .QN(n19342) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n3132), .CK(CLK), .RN(n19056), .QN(
        n19632) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n3131), .CK(CLK), .RN(n19056), .QN(
        n19633) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n3130), .CK(CLK), .RN(n19056), .QN(
        n19634) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n3129), .CK(CLK), .RN(n19056), .QN(
        n19635) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n3128), .CK(CLK), .RN(n19056), .QN(
        n19636) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n3127), .CK(CLK), .RN(n19056), .QN(
        n19637) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n3126), .CK(CLK), .RN(n19056), .QN(
        n19638) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n3125), .CK(CLK), .RN(n19056), .QN(
        n19751) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n3124), .CK(CLK), .RN(n19056), .QN(
        n19752) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n3123), .CK(CLK), .RN(n19056), .QN(
        n19753) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n3122), .CK(CLK), .RN(n19056), .QN(
        n19754) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n3121), .CK(CLK), .RN(n19056), .QN(
        n19755) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n3120), .CK(CLK), .RN(n19056), .QN(
        n19756) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n3119), .CK(CLK), .RN(n19056), .QN(
        n19757) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n3118), .CK(CLK), .RN(n19056), .QN(
        n19758) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n3117), .CK(CLK), .RN(n19056), .QN(
        n19759) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n3116), .CK(CLK), .RN(n19056), .QN(
        n19760) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n3115), .CK(CLK), .RN(n19056), .QN(
        n19761) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n3114), .CK(CLK), .RN(n19056), .QN(
        n19762) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n3113), .CK(CLK), .RN(n19056), .QN(
        n19763) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n3112), .CK(CLK), .RN(n19056), .QN(
        n19764) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n3104), .CK(CLK), .RN(n19056), .QN(
        n19772) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n3103), .CK(CLK), .RN(n19056), .QN(
        n19773) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n3102), .CK(CLK), .RN(n19056), .QN(
        n19774) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n3260), .CK(CLK), .RN(n19056), .Q(
        n17669), .QN(n19648) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n3259), .CK(CLK), .RN(n19056), .Q(
        n17668), .QN(n19649) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n3258), .CK(CLK), .RN(n19056), .Q(
        n17667), .QN(n19650) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n3257), .CK(CLK), .RN(n19056), .Q(
        n17666), .QN(n19651) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n3256), .CK(CLK), .RN(n19056), .Q(
        n17665), .QN(n19652) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n3255), .CK(CLK), .RN(n19056), .Q(
        n17664), .QN(n19653) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n3254), .CK(CLK), .RN(n19056), .Q(
        n17663), .QN(n19654) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n3253), .CK(CLK), .RN(n19056), .Q(
        n17550), .QN(n19799) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n3252), .CK(CLK), .RN(n19056), .Q(
        n17549), .QN(n19800) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n3251), .CK(CLK), .RN(n19056), .Q(
        n17548), .QN(n19801) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n3250), .CK(CLK), .RN(n19056), .Q(
        n17547), .QN(n19802) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n3249), .CK(CLK), .RN(n19056), .Q(
        n17546), .QN(n19803) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n3248), .CK(CLK), .RN(n19056), .Q(
        n17545), .QN(n19804) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n3247), .CK(CLK), .RN(n19056), .Q(
        n17544), .QN(n19805) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n3246), .CK(CLK), .RN(n19056), .Q(
        n17543), .QN(n19806) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n3245), .CK(CLK), .RN(n19056), .Q(
        n17542), .QN(n19807) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n3244), .CK(CLK), .RN(n19056), .Q(
        n17541), .QN(n19808) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n3243), .CK(CLK), .RN(n19056), .Q(
        n17540), .QN(n19809) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n3242), .CK(CLK), .RN(n19056), .Q(
        n17539), .QN(n19810) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n3241), .CK(CLK), .RN(n19056), .Q(
        n17538), .QN(n19811) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n3240), .CK(CLK), .RN(n19056), .Q(
        n17537), .QN(n19812) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n3232), .CK(CLK), .RN(n19056), .Q(n17529), .QN(n19820) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n3231), .CK(CLK), .RN(n19056), .Q(n17528), .QN(n19821) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n3230), .CK(CLK), .RN(n19056), .Q(n17527), .QN(n19822) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n3292), .CK(CLK), .RN(n19056), .Q(
        n17685), .QN(n19616) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n3291), .CK(CLK), .RN(n19056), .Q(
        n17684), .QN(n19617) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n3290), .CK(CLK), .RN(n19056), .Q(
        n17683), .QN(n19618) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n3289), .CK(CLK), .RN(n19056), .Q(
        n17682), .QN(n19619) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n3288), .CK(CLK), .RN(n19056), .Q(
        n17681), .QN(n19620) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n3287), .CK(CLK), .RN(n19056), .Q(
        n17680), .QN(n19621) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n3286), .CK(CLK), .RN(n19056), .Q(
        n17679), .QN(n19622) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n3285), .CK(CLK), .RN(n19056), .Q(
        n17598), .QN(n19703) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n3284), .CK(CLK), .RN(n19056), .Q(
        n17597), .QN(n19704) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n3283), .CK(CLK), .RN(n19056), .Q(
        n17596), .QN(n19705) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n3282), .CK(CLK), .RN(n19056), .Q(
        n17595), .QN(n19706) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n3281), .CK(CLK), .RN(n19056), .Q(
        n17594), .QN(n19707) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n3280), .CK(CLK), .RN(n19056), .Q(
        n17593), .QN(n19708) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n3279), .CK(CLK), .RN(n19056), .Q(
        n17592), .QN(n19709) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n3278), .CK(CLK), .RN(n19056), .Q(
        n17591), .QN(n19710) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n3277), .CK(CLK), .RN(n19056), .Q(
        n17590), .QN(n19711) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n3276), .CK(CLK), .RN(n19056), .Q(
        n17589), .QN(n19712) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n3275), .CK(CLK), .RN(n19056), .Q(
        n17588), .QN(n19713) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n3274), .CK(CLK), .RN(n19056), .Q(
        n17587), .QN(n19714) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n3273), .CK(CLK), .RN(n19056), .Q(
        n17586), .QN(n19715) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n3272), .CK(CLK), .RN(n19056), .Q(
        n17585), .QN(n19716) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n3264), .CK(CLK), .RN(n19056), .Q(n17577), .QN(n19724) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n3263), .CK(CLK), .RN(n19056), .Q(n17576), .QN(n19725) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n3262), .CK(CLK), .RN(n19056), .Q(n17575), .QN(n19726) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n3388), .CK(CLK), .RN(n19056), .QN(
        n19656) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n3387), .CK(CLK), .RN(n19056), .QN(
        n19657) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n3386), .CK(CLK), .RN(n19056), .QN(
        n19658) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n3385), .CK(CLK), .RN(n19056), .QN(
        n19659) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n3384), .CK(CLK), .RN(n19056), .QN(
        n19660) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n3383), .CK(CLK), .RN(n19056), .QN(
        n19661) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n3382), .CK(CLK), .RN(n19056), .QN(
        n19662) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n3360), .CK(CLK), .RN(n19056), .QN(n19830) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n3359), .CK(CLK), .RN(n19056), .QN(n19831) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n3358), .CK(CLK), .RN(n19056), .QN(n19832) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n19059), .CK(CLK), .RN(n19056), .Q(
        n17622) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n19061), .CK(CLK), .RN(n19056), .Q(
        n17621) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n19063), .CK(CLK), .RN(n19056), .Q(
        n17620) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n19065), .CK(CLK), .RN(n19056), .Q(
        n17619) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n19067), .CK(CLK), .RN(n19056), .Q(
        n17618) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n19069), .CK(CLK), .RN(n19056), .Q(
        n17617) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n19071), .CK(CLK), .RN(n19056), .Q(
        n17616) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n19073), .CK(CLK), .RN(n19056), .Q(
        n17615) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n19075), .CK(CLK), .RN(n19056), .Q(
        n17614) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n19077), .CK(CLK), .RN(n19056), .Q(
        n17613) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n19079), .CK(CLK), .RN(n19056), .Q(
        n17612) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n19081), .CK(CLK), .RN(n19056), .Q(
        n17611) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n19083), .CK(CLK), .RN(n19056), .Q(
        n17610) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n19085), .CK(CLK), .RN(n19056), .Q(
        n17609) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n19087), .CK(CLK), .RN(n19056), .Q(
        n17608) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n19089), .CK(CLK), .RN(n19056), .Q(
        n17607) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n19091), .CK(CLK), .RN(n19056), .Q(
        n17606) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n19093), .CK(CLK), .RN(n19056), .Q(
        n17605) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n19095), .CK(CLK), .RN(n19056), .Q(
        n17604) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n19097), .CK(CLK), .RN(n19056), .Q(
        n17603) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n19099), .CK(CLK), .RN(n19056), .Q(
        n17602) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n19101), .CK(CLK), .RN(n19056), .Q(
        n17601) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n19103), .CK(CLK), .RN(n19056), .Q(
        n17600) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n19105), .CK(CLK), .RN(n19056), .Q(
        n17599) );
  INV_X1 U2 ( .A(ADD_RD1[2]), .ZN(n19913) );
  AND3_X1 U3 ( .A1(ADD_RD1[3]), .A2(n19915), .A3(RD1), .ZN(n1583) );
  AND3_X1 U4 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .A3(RD1), .ZN(n1573) );
  AND3_X1 U5 ( .A1(ADD_RD1[4]), .A2(n19916), .A3(RD1), .ZN(n1574) );
  AND2_X1 U6 ( .A1(n937), .A2(n899), .ZN(n18389) );
  AND2_X1 U7 ( .A1(n902), .A2(n899), .ZN(n18390) );
  AND2_X1 U8 ( .A1(n940), .A2(n899), .ZN(n18391) );
  AND2_X1 U9 ( .A1(n940), .A2(n936), .ZN(n18392) );
  AND2_X1 U10 ( .A1(n957), .A2(n939), .ZN(n18393) );
  AND2_X1 U11 ( .A1(n957), .A2(n899), .ZN(n18394) );
  AND2_X1 U12 ( .A1(n954), .A2(n936), .ZN(n18395) );
  AND2_X1 U13 ( .A1(n959), .A2(n939), .ZN(n18396) );
  AND2_X1 U14 ( .A1(n959), .A2(n943), .ZN(n18397) );
  AND2_X1 U15 ( .A1(n959), .A2(n899), .ZN(n18398) );
  AND2_X1 U16 ( .A1(n961), .A2(n943), .ZN(n18399) );
  AND2_X1 U17 ( .A1(n961), .A2(n899), .ZN(n18400) );
  AND2_X1 U18 ( .A1(n954), .A2(n943), .ZN(n18401) );
  AND2_X1 U19 ( .A1(n957), .A2(n943), .ZN(n18402) );
  AND2_X1 U20 ( .A1(n961), .A2(n939), .ZN(n18403) );
  AND2_X1 U21 ( .A1(n961), .A2(n936), .ZN(n18404) );
  AND2_X1 U22 ( .A1(n954), .A2(n899), .ZN(n18405) );
  AND2_X1 U23 ( .A1(n959), .A2(n936), .ZN(n18406) );
  AND2_X1 U24 ( .A1(n954), .A2(n939), .ZN(n18407) );
  AND2_X1 U25 ( .A1(n957), .A2(n936), .ZN(n18408) );
  AND2_X1 U26 ( .A1(n939), .A2(n937), .ZN(n18409) );
  AND2_X1 U27 ( .A1(n939), .A2(n902), .ZN(n18410) );
  AND2_X1 U28 ( .A1(n936), .A2(n902), .ZN(n18411) );
  AND2_X1 U29 ( .A1(n943), .A2(n900), .ZN(n18412) );
  AND2_X1 U30 ( .A1(n939), .A2(n900), .ZN(n18413) );
  AND2_X1 U31 ( .A1(n943), .A2(n902), .ZN(n18414) );
  AND2_X1 U32 ( .A1(n936), .A2(n900), .ZN(n18415) );
  AND2_X1 U33 ( .A1(n943), .A2(n937), .ZN(n18416) );
  AND2_X1 U34 ( .A1(n943), .A2(n940), .ZN(n18417) );
  AND2_X1 U35 ( .A1(n939), .A2(n940), .ZN(n18418) );
  INV_X32 U36 ( .A(n19055), .ZN(n19056) );
  CLKBUF_X1 U37 ( .A(RESET), .Z(n19055) );
  INV_X1 U38 ( .A(n18849), .ZN(n18839) );
  INV_X1 U39 ( .A(n18849), .ZN(n18840) );
  INV_X1 U40 ( .A(n18728), .ZN(n18719) );
  INV_X1 U41 ( .A(n18728), .ZN(n18718) );
  INV_X1 U42 ( .A(n18948), .ZN(n18939) );
  INV_X1 U43 ( .A(n18948), .ZN(n18938) );
  INV_X1 U44 ( .A(n18992), .ZN(n18983) );
  INV_X1 U45 ( .A(n18992), .ZN(n18982) );
  INV_X1 U46 ( .A(n18827), .ZN(n18817) );
  INV_X1 U47 ( .A(n18827), .ZN(n18818) );
  INV_X1 U48 ( .A(n18937), .ZN(n18928) );
  INV_X1 U49 ( .A(n18937), .ZN(n18927) );
  INV_X1 U50 ( .A(n18783), .ZN(n18773) );
  INV_X1 U51 ( .A(n18783), .ZN(n18774) );
  INV_X1 U52 ( .A(n18970), .ZN(n18961) );
  INV_X1 U53 ( .A(n18970), .ZN(n18960) );
  INV_X1 U54 ( .A(n18838), .ZN(n18828) );
  INV_X1 U55 ( .A(n18838), .ZN(n18829) );
  INV_X1 U56 ( .A(n18904), .ZN(n18895) );
  INV_X1 U57 ( .A(n18904), .ZN(n18894) );
  INV_X1 U58 ( .A(n19014), .ZN(n19004) );
  INV_X1 U59 ( .A(n19014), .ZN(n19005) );
  INV_X1 U60 ( .A(n18959), .ZN(n18950) );
  INV_X1 U61 ( .A(n18959), .ZN(n18949) );
  INV_X1 U62 ( .A(n18794), .ZN(n18784) );
  INV_X1 U63 ( .A(n18794), .ZN(n18785) );
  INV_X1 U64 ( .A(n18761), .ZN(n18751) );
  INV_X1 U65 ( .A(n18761), .ZN(n18752) );
  INV_X1 U66 ( .A(n18860), .ZN(n18850) );
  INV_X1 U67 ( .A(n18860), .ZN(n18851) );
  INV_X1 U68 ( .A(n18816), .ZN(n18806) );
  INV_X1 U69 ( .A(n18816), .ZN(n18807) );
  INV_X1 U70 ( .A(n18772), .ZN(n18762) );
  INV_X1 U71 ( .A(n18772), .ZN(n18763) );
  INV_X1 U72 ( .A(n18739), .ZN(n18729) );
  INV_X1 U73 ( .A(n18739), .ZN(n18730) );
  INV_X1 U74 ( .A(n18893), .ZN(n18884) );
  INV_X1 U75 ( .A(n18893), .ZN(n18883) );
  INV_X1 U76 ( .A(n18871), .ZN(n18861) );
  INV_X1 U77 ( .A(n18871), .ZN(n18862) );
  INV_X1 U78 ( .A(n18915), .ZN(n18906) );
  INV_X1 U79 ( .A(n18915), .ZN(n18905) );
  INV_X1 U80 ( .A(n18750), .ZN(n18740) );
  INV_X1 U81 ( .A(n18750), .ZN(n18741) );
  INV_X1 U82 ( .A(n19003), .ZN(n18993) );
  INV_X1 U83 ( .A(n19003), .ZN(n18994) );
  INV_X1 U84 ( .A(n18926), .ZN(n18917) );
  INV_X1 U85 ( .A(n18926), .ZN(n18916) );
  INV_X1 U86 ( .A(n18981), .ZN(n18972) );
  INV_X1 U87 ( .A(n18981), .ZN(n18971) );
  INV_X1 U88 ( .A(n18882), .ZN(n18872) );
  INV_X1 U89 ( .A(n18882), .ZN(n18873) );
  INV_X1 U90 ( .A(n19025), .ZN(n19015) );
  INV_X1 U91 ( .A(n19025), .ZN(n19016) );
  INV_X1 U92 ( .A(n18805), .ZN(n18795) );
  INV_X1 U93 ( .A(n18805), .ZN(n18796) );
  INV_X1 U94 ( .A(n19045), .ZN(n19035) );
  INV_X1 U95 ( .A(n19045), .ZN(n19036) );
  INV_X1 U96 ( .A(n18717), .ZN(n18708) );
  INV_X1 U97 ( .A(n18717), .ZN(n18707) );
  BUF_X1 U98 ( .A(n18399), .Z(n18849) );
  BUF_X1 U99 ( .A(n18843), .Z(n18848) );
  BUF_X1 U100 ( .A(n18842), .Z(n18847) );
  BUF_X1 U101 ( .A(n18399), .Z(n18846) );
  BUF_X1 U102 ( .A(n18399), .Z(n18845) );
  BUF_X1 U103 ( .A(n18399), .Z(n18844) );
  BUF_X1 U104 ( .A(n18399), .Z(n18843) );
  BUF_X1 U105 ( .A(n18399), .Z(n18842) );
  BUF_X1 U106 ( .A(n18399), .Z(n18841) );
  INV_X1 U107 ( .A(n19034), .ZN(n19027) );
  INV_X1 U108 ( .A(n19034), .ZN(n19026) );
  INV_X1 U109 ( .A(n19054), .ZN(n19046) );
  INV_X1 U110 ( .A(n19054), .ZN(n19047) );
  BUF_X1 U111 ( .A(n18390), .Z(n19045) );
  BUF_X1 U112 ( .A(n18404), .Z(n18728) );
  BUF_X1 U113 ( .A(n18391), .Z(n18948) );
  BUF_X1 U114 ( .A(n18392), .Z(n18992) );
  BUF_X1 U115 ( .A(n18389), .Z(n18794) );
  BUF_X1 U116 ( .A(n18393), .Z(n18827) );
  BUF_X1 U117 ( .A(n18405), .Z(n18937) );
  BUF_X1 U118 ( .A(n18394), .Z(n18783) );
  BUF_X1 U119 ( .A(n18395), .Z(n18970) );
  BUF_X1 U120 ( .A(n18402), .Z(n18871) );
  BUF_X1 U121 ( .A(n18400), .Z(n18761) );
  BUF_X1 U122 ( .A(n18397), .Z(n18860) );
  BUF_X1 U123 ( .A(n18396), .Z(n18816) );
  BUF_X1 U124 ( .A(n18398), .Z(n18772) );
  BUF_X1 U125 ( .A(n18406), .Z(n18739) );
  BUF_X1 U126 ( .A(n18401), .Z(n18893) );
  BUF_X1 U127 ( .A(n18407), .Z(n18915) );
  BUF_X1 U128 ( .A(n18408), .Z(n18750) );
  BUF_X1 U129 ( .A(n18403), .Z(n18805) );
  BUF_X1 U130 ( .A(n18409), .Z(n18838) );
  BUF_X1 U131 ( .A(n18417), .Z(n18904) );
  BUF_X1 U132 ( .A(n18410), .Z(n19014) );
  BUF_X1 U133 ( .A(n18411), .Z(n18959) );
  BUF_X1 U134 ( .A(n18412), .Z(n19003) );
  BUF_X1 U135 ( .A(n18413), .Z(n18926) );
  BUF_X1 U136 ( .A(n18415), .Z(n18981) );
  BUF_X1 U137 ( .A(n18416), .Z(n18882) );
  BUF_X1 U138 ( .A(n18418), .Z(n19025) );
  BUF_X1 U139 ( .A(n18414), .Z(n18717) );
  BUF_X1 U140 ( .A(n18788), .Z(n18793) );
  BUF_X1 U141 ( .A(n18787), .Z(n18792) );
  BUF_X1 U142 ( .A(n18389), .Z(n18791) );
  BUF_X1 U143 ( .A(n18389), .Z(n18790) );
  BUF_X1 U144 ( .A(n18389), .Z(n18789) );
  BUF_X1 U145 ( .A(n18389), .Z(n18788) );
  BUF_X1 U146 ( .A(n18389), .Z(n18787) );
  BUF_X1 U147 ( .A(n18389), .Z(n18786) );
  BUF_X1 U148 ( .A(n19039), .Z(n19044) );
  BUF_X1 U149 ( .A(n19038), .Z(n19043) );
  BUF_X1 U150 ( .A(n18390), .Z(n19042) );
  BUF_X1 U151 ( .A(n18390), .Z(n19041) );
  BUF_X1 U152 ( .A(n18390), .Z(n19040) );
  BUF_X1 U153 ( .A(n18390), .Z(n19039) );
  BUF_X1 U154 ( .A(n18390), .Z(n19038) );
  BUF_X1 U155 ( .A(n18390), .Z(n19037) );
  BUF_X1 U156 ( .A(n18404), .Z(n18720) );
  BUF_X1 U157 ( .A(n18404), .Z(n18721) );
  BUF_X1 U158 ( .A(n18404), .Z(n18722) );
  BUF_X1 U159 ( .A(n18404), .Z(n18723) );
  BUF_X1 U160 ( .A(n18404), .Z(n18724) );
  BUF_X1 U161 ( .A(n18404), .Z(n18725) );
  BUF_X1 U162 ( .A(n18723), .Z(n18726) );
  BUF_X1 U163 ( .A(n18724), .Z(n18727) );
  BUF_X1 U164 ( .A(n18405), .Z(n18931) );
  BUF_X1 U165 ( .A(n18405), .Z(n18932) );
  BUF_X1 U166 ( .A(n18405), .Z(n18933) );
  BUF_X1 U167 ( .A(n18405), .Z(n18934) );
  BUF_X1 U168 ( .A(n18931), .Z(n18935) );
  BUF_X1 U169 ( .A(n18929), .Z(n18936) );
  BUF_X1 U170 ( .A(n18405), .Z(n18929) );
  BUF_X1 U171 ( .A(n18405), .Z(n18930) );
  BUF_X1 U172 ( .A(n18756), .Z(n18760) );
  BUF_X1 U173 ( .A(n18755), .Z(n18759) );
  BUF_X1 U174 ( .A(n18400), .Z(n18758) );
  BUF_X1 U175 ( .A(n18400), .Z(n18757) );
  BUF_X1 U176 ( .A(n18400), .Z(n18756) );
  BUF_X1 U177 ( .A(n18400), .Z(n18755) );
  BUF_X1 U178 ( .A(n18854), .Z(n18859) );
  BUF_X1 U179 ( .A(n18853), .Z(n18858) );
  BUF_X1 U180 ( .A(n18397), .Z(n18857) );
  BUF_X1 U181 ( .A(n18397), .Z(n18856) );
  BUF_X1 U182 ( .A(n18397), .Z(n18855) );
  BUF_X1 U183 ( .A(n18397), .Z(n18854) );
  BUF_X1 U184 ( .A(n18810), .Z(n18815) );
  BUF_X1 U185 ( .A(n18809), .Z(n18814) );
  BUF_X1 U186 ( .A(n18396), .Z(n18813) );
  BUF_X1 U187 ( .A(n18396), .Z(n18812) );
  BUF_X1 U188 ( .A(n18396), .Z(n18811) );
  BUF_X1 U189 ( .A(n18396), .Z(n18810) );
  BUF_X1 U190 ( .A(n18766), .Z(n18771) );
  BUF_X1 U191 ( .A(n18765), .Z(n18770) );
  BUF_X1 U192 ( .A(n18398), .Z(n18769) );
  BUF_X1 U193 ( .A(n18398), .Z(n18768) );
  BUF_X1 U194 ( .A(n18398), .Z(n18767) );
  BUF_X1 U195 ( .A(n18398), .Z(n18766) );
  BUF_X1 U196 ( .A(n18733), .Z(n18737) );
  BUF_X1 U197 ( .A(n18406), .Z(n18736) );
  BUF_X1 U198 ( .A(n18406), .Z(n18735) );
  BUF_X1 U199 ( .A(n18406), .Z(n18734) );
  BUF_X1 U200 ( .A(n18736), .Z(n18738) );
  BUF_X1 U201 ( .A(n18406), .Z(n18733) );
  BUF_X1 U202 ( .A(n18401), .Z(n18887) );
  BUF_X1 U203 ( .A(n18401), .Z(n18888) );
  BUF_X1 U204 ( .A(n18401), .Z(n18889) );
  BUF_X1 U205 ( .A(n18401), .Z(n18890) );
  BUF_X1 U206 ( .A(n18887), .Z(n18891) );
  BUF_X1 U207 ( .A(n18885), .Z(n18892) );
  BUF_X1 U208 ( .A(n18402), .Z(n18865) );
  BUF_X1 U209 ( .A(n18402), .Z(n18864) );
  BUF_X1 U210 ( .A(n18402), .Z(n18863) );
  BUF_X1 U211 ( .A(n18407), .Z(n18909) );
  BUF_X1 U212 ( .A(n18407), .Z(n18910) );
  BUF_X1 U213 ( .A(n18407), .Z(n18911) );
  BUF_X1 U214 ( .A(n18407), .Z(n18912) );
  BUF_X1 U215 ( .A(n18909), .Z(n18913) );
  BUF_X1 U216 ( .A(n18907), .Z(n18914) );
  BUF_X1 U217 ( .A(n18744), .Z(n18749) );
  BUF_X1 U218 ( .A(n18747), .Z(n18748) );
  BUF_X1 U219 ( .A(n18408), .Z(n18747) );
  BUF_X1 U220 ( .A(n18408), .Z(n18746) );
  BUF_X1 U221 ( .A(n18408), .Z(n18745) );
  BUF_X1 U222 ( .A(n18408), .Z(n18744) );
  BUF_X1 U223 ( .A(n18799), .Z(n18804) );
  BUF_X1 U224 ( .A(n18798), .Z(n18803) );
  BUF_X1 U225 ( .A(n18403), .Z(n18802) );
  BUF_X1 U226 ( .A(n18403), .Z(n18801) );
  BUF_X1 U227 ( .A(n18403), .Z(n18800) );
  BUF_X1 U228 ( .A(n18403), .Z(n18799) );
  BUF_X1 U229 ( .A(n18400), .Z(n18754) );
  BUF_X1 U230 ( .A(n18400), .Z(n18753) );
  BUF_X1 U231 ( .A(n18397), .Z(n18853) );
  BUF_X1 U232 ( .A(n18397), .Z(n18852) );
  BUF_X1 U233 ( .A(n18396), .Z(n18809) );
  BUF_X1 U234 ( .A(n18396), .Z(n18808) );
  BUF_X1 U235 ( .A(n18398), .Z(n18765) );
  BUF_X1 U236 ( .A(n18398), .Z(n18764) );
  BUF_X1 U237 ( .A(n18406), .Z(n18732) );
  BUF_X1 U238 ( .A(n18406), .Z(n18731) );
  BUF_X1 U239 ( .A(n18401), .Z(n18885) );
  BUF_X1 U240 ( .A(n18401), .Z(n18886) );
  BUF_X1 U241 ( .A(n18407), .Z(n18907) );
  BUF_X1 U242 ( .A(n18407), .Z(n18908) );
  BUF_X1 U243 ( .A(n18408), .Z(n18743) );
  BUF_X1 U244 ( .A(n18408), .Z(n18742) );
  BUF_X1 U245 ( .A(n18403), .Z(n18798) );
  BUF_X1 U246 ( .A(n18403), .Z(n18797) );
  BUF_X1 U247 ( .A(n18417), .Z(n18898) );
  BUF_X1 U248 ( .A(n18417), .Z(n18899) );
  BUF_X1 U249 ( .A(n18417), .Z(n18900) );
  BUF_X1 U250 ( .A(n18417), .Z(n18901) );
  BUF_X1 U251 ( .A(n18898), .Z(n18902) );
  BUF_X1 U252 ( .A(n18896), .Z(n18903) );
  BUF_X1 U253 ( .A(n18417), .Z(n18896) );
  BUF_X1 U254 ( .A(n18417), .Z(n18897) );
  BUF_X1 U255 ( .A(n18412), .Z(n18995) );
  BUF_X1 U256 ( .A(n18415), .Z(n18975) );
  BUF_X1 U257 ( .A(n18415), .Z(n18976) );
  BUF_X1 U258 ( .A(n18415), .Z(n18977) );
  BUF_X1 U259 ( .A(n18415), .Z(n18978) );
  BUF_X1 U260 ( .A(n18975), .Z(n18979) );
  BUF_X1 U261 ( .A(n18973), .Z(n18980) );
  BUF_X1 U262 ( .A(n18876), .Z(n18881) );
  BUF_X1 U263 ( .A(n18875), .Z(n18880) );
  BUF_X1 U264 ( .A(n18416), .Z(n18879) );
  BUF_X1 U265 ( .A(n18416), .Z(n18878) );
  BUF_X1 U266 ( .A(n18416), .Z(n18877) );
  BUF_X1 U267 ( .A(n18416), .Z(n18876) );
  BUF_X1 U268 ( .A(n19019), .Z(n19024) );
  BUF_X1 U269 ( .A(n19018), .Z(n19023) );
  BUF_X1 U270 ( .A(n18418), .Z(n19022) );
  BUF_X1 U271 ( .A(n18418), .Z(n19021) );
  BUF_X1 U272 ( .A(n18418), .Z(n19020) );
  BUF_X1 U273 ( .A(n18418), .Z(n19019) );
  BUF_X1 U274 ( .A(n18415), .Z(n18973) );
  BUF_X1 U275 ( .A(n18415), .Z(n18974) );
  BUF_X1 U276 ( .A(n18416), .Z(n18875) );
  BUF_X1 U277 ( .A(n18416), .Z(n18874) );
  BUF_X1 U278 ( .A(n18418), .Z(n19018) );
  BUF_X1 U279 ( .A(n18418), .Z(n19017) );
  BUF_X1 U280 ( .A(n18402), .Z(n18866) );
  BUF_X1 U281 ( .A(n18413), .Z(n18918) );
  BUF_X1 U282 ( .A(n18391), .Z(n18942) );
  BUF_X1 U283 ( .A(n18391), .Z(n18943) );
  BUF_X1 U284 ( .A(n18391), .Z(n18944) );
  BUF_X1 U285 ( .A(n18391), .Z(n18945) );
  BUF_X1 U286 ( .A(n18942), .Z(n18946) );
  BUF_X1 U287 ( .A(n18940), .Z(n18947) );
  BUF_X1 U288 ( .A(n18392), .Z(n18986) );
  BUF_X1 U289 ( .A(n18392), .Z(n18987) );
  BUF_X1 U290 ( .A(n18392), .Z(n18988) );
  BUF_X1 U291 ( .A(n18392), .Z(n18989) );
  BUF_X1 U292 ( .A(n18986), .Z(n18990) );
  BUF_X1 U293 ( .A(n18984), .Z(n18991) );
  BUF_X1 U294 ( .A(n18865), .Z(n18870) );
  BUF_X1 U295 ( .A(n18864), .Z(n18869) );
  BUF_X1 U296 ( .A(n18821), .Z(n18826) );
  BUF_X1 U297 ( .A(n18820), .Z(n18825) );
  BUF_X1 U298 ( .A(n18393), .Z(n18824) );
  BUF_X1 U299 ( .A(n18393), .Z(n18823) );
  BUF_X1 U300 ( .A(n18393), .Z(n18822) );
  BUF_X1 U301 ( .A(n18393), .Z(n18821) );
  BUF_X1 U302 ( .A(n18777), .Z(n18782) );
  BUF_X1 U303 ( .A(n18776), .Z(n18781) );
  BUF_X1 U304 ( .A(n18394), .Z(n18780) );
  BUF_X1 U305 ( .A(n18394), .Z(n18779) );
  BUF_X1 U306 ( .A(n18394), .Z(n18778) );
  BUF_X1 U307 ( .A(n18394), .Z(n18777) );
  BUF_X1 U308 ( .A(n18395), .Z(n18964) );
  BUF_X1 U309 ( .A(n18395), .Z(n18965) );
  BUF_X1 U310 ( .A(n18395), .Z(n18966) );
  BUF_X1 U311 ( .A(n18395), .Z(n18967) );
  BUF_X1 U312 ( .A(n18964), .Z(n18968) );
  BUF_X1 U313 ( .A(n18962), .Z(n18969) );
  BUF_X1 U314 ( .A(n18391), .Z(n18940) );
  BUF_X1 U315 ( .A(n18391), .Z(n18941) );
  BUF_X1 U316 ( .A(n18392), .Z(n18984) );
  BUF_X1 U317 ( .A(n18392), .Z(n18985) );
  BUF_X1 U318 ( .A(n18402), .Z(n18867) );
  BUF_X1 U319 ( .A(n18402), .Z(n18868) );
  BUF_X1 U320 ( .A(n18393), .Z(n18820) );
  BUF_X1 U321 ( .A(n18393), .Z(n18819) );
  BUF_X1 U322 ( .A(n18394), .Z(n18776) );
  BUF_X1 U323 ( .A(n18394), .Z(n18775) );
  BUF_X1 U324 ( .A(n18395), .Z(n18962) );
  BUF_X1 U325 ( .A(n18395), .Z(n18963) );
  BUF_X1 U326 ( .A(n18832), .Z(n18837) );
  BUF_X1 U327 ( .A(n18831), .Z(n18836) );
  BUF_X1 U328 ( .A(n18409), .Z(n18835) );
  BUF_X1 U329 ( .A(n18409), .Z(n18834) );
  BUF_X1 U330 ( .A(n18409), .Z(n18833) );
  BUF_X1 U331 ( .A(n18409), .Z(n18832) );
  BUF_X1 U332 ( .A(n18409), .Z(n18831) );
  BUF_X1 U333 ( .A(n18409), .Z(n18830) );
  BUF_X1 U334 ( .A(n19008), .Z(n19013) );
  BUF_X1 U335 ( .A(n19007), .Z(n19012) );
  BUF_X1 U336 ( .A(n18410), .Z(n19011) );
  BUF_X1 U337 ( .A(n18410), .Z(n19010) );
  BUF_X1 U338 ( .A(n18410), .Z(n19009) );
  BUF_X1 U339 ( .A(n18410), .Z(n19008) );
  BUF_X1 U340 ( .A(n18411), .Z(n18953) );
  BUF_X1 U341 ( .A(n18411), .Z(n18954) );
  BUF_X1 U342 ( .A(n18411), .Z(n18955) );
  BUF_X1 U343 ( .A(n18411), .Z(n18956) );
  BUF_X1 U344 ( .A(n18953), .Z(n18957) );
  BUF_X1 U345 ( .A(n18951), .Z(n18958) );
  BUF_X1 U346 ( .A(n18410), .Z(n19007) );
  BUF_X1 U347 ( .A(n18410), .Z(n19006) );
  BUF_X1 U348 ( .A(n18411), .Z(n18951) );
  BUF_X1 U349 ( .A(n18411), .Z(n18952) );
  BUF_X1 U350 ( .A(n18995), .Z(n19002) );
  BUF_X1 U351 ( .A(n18997), .Z(n19001) );
  BUF_X1 U352 ( .A(n18412), .Z(n19000) );
  BUF_X1 U353 ( .A(n18413), .Z(n18920) );
  BUF_X1 U354 ( .A(n18413), .Z(n18921) );
  BUF_X1 U355 ( .A(n18413), .Z(n18923) );
  BUF_X1 U356 ( .A(n18918), .Z(n18924) );
  BUF_X1 U357 ( .A(n18920), .Z(n18925) );
  BUF_X1 U358 ( .A(n18412), .Z(n18998) );
  BUF_X1 U359 ( .A(n18412), .Z(n18997) );
  BUF_X1 U360 ( .A(n18412), .Z(n18996) );
  BUF_X1 U361 ( .A(n18412), .Z(n18999) );
  BUF_X1 U362 ( .A(n18413), .Z(n18922) );
  BUF_X1 U363 ( .A(n18413), .Z(n18919) );
  BUF_X1 U364 ( .A(n18414), .Z(n18711) );
  BUF_X1 U365 ( .A(n18414), .Z(n18712) );
  BUF_X1 U366 ( .A(n18414), .Z(n18713) );
  BUF_X1 U367 ( .A(n18414), .Z(n18714) );
  BUF_X1 U368 ( .A(n18711), .Z(n18715) );
  BUF_X1 U369 ( .A(n18712), .Z(n18716) );
  BUF_X1 U370 ( .A(n18414), .Z(n18709) );
  BUF_X1 U371 ( .A(n18414), .Z(n18710) );
  BUF_X1 U372 ( .A(n19120), .Z(n18512) );
  BUF_X1 U373 ( .A(n19118), .Z(n18509) );
  BUF_X1 U374 ( .A(n19116), .Z(n18506) );
  BUF_X1 U375 ( .A(n19114), .Z(n18503) );
  BUF_X1 U376 ( .A(n19112), .Z(n18500) );
  BUF_X1 U377 ( .A(n19110), .Z(n18497) );
  BUF_X1 U378 ( .A(n19108), .Z(n18494) );
  BUF_X1 U379 ( .A(n19106), .Z(n18491) );
  BUF_X1 U380 ( .A(n19104), .Z(n18488) );
  BUF_X1 U381 ( .A(n19102), .Z(n18485) );
  BUF_X1 U382 ( .A(n19100), .Z(n18482) );
  BUF_X1 U383 ( .A(n19098), .Z(n18479) );
  BUF_X1 U384 ( .A(n19096), .Z(n18476) );
  BUF_X1 U385 ( .A(n19094), .Z(n18473) );
  BUF_X1 U386 ( .A(n19092), .Z(n18470) );
  BUF_X1 U387 ( .A(n19090), .Z(n18467) );
  BUF_X1 U388 ( .A(n19088), .Z(n18464) );
  BUF_X1 U389 ( .A(n19086), .Z(n18461) );
  BUF_X1 U390 ( .A(n19084), .Z(n18458) );
  BUF_X1 U391 ( .A(n19082), .Z(n18455) );
  BUF_X1 U392 ( .A(n19080), .Z(n18452) );
  BUF_X1 U393 ( .A(n19078), .Z(n18449) );
  BUF_X1 U394 ( .A(n19076), .Z(n18446) );
  BUF_X1 U395 ( .A(n19074), .Z(n18443) );
  BUF_X1 U396 ( .A(n19072), .Z(n18440) );
  BUF_X1 U397 ( .A(n19070), .Z(n18437) );
  BUF_X1 U398 ( .A(n19068), .Z(n18434) );
  BUF_X1 U399 ( .A(n19066), .Z(n18431) );
  BUF_X1 U400 ( .A(n19064), .Z(n18428) );
  BUF_X1 U401 ( .A(n19062), .Z(n18425) );
  BUF_X1 U402 ( .A(n19060), .Z(n18422) );
  BUF_X1 U403 ( .A(n19058), .Z(n18419) );
  BUF_X1 U404 ( .A(n19104), .Z(n18489) );
  BUF_X1 U405 ( .A(n19102), .Z(n18486) );
  BUF_X1 U406 ( .A(n19100), .Z(n18483) );
  BUF_X1 U407 ( .A(n19098), .Z(n18480) );
  BUF_X1 U408 ( .A(n19096), .Z(n18477) );
  BUF_X1 U409 ( .A(n19094), .Z(n18474) );
  BUF_X1 U410 ( .A(n19092), .Z(n18471) );
  BUF_X1 U411 ( .A(n19090), .Z(n18468) );
  BUF_X1 U412 ( .A(n19088), .Z(n18465) );
  BUF_X1 U413 ( .A(n19086), .Z(n18462) );
  BUF_X1 U414 ( .A(n19084), .Z(n18459) );
  BUF_X1 U415 ( .A(n19082), .Z(n18456) );
  BUF_X1 U416 ( .A(n19080), .Z(n18453) );
  BUF_X1 U417 ( .A(n19078), .Z(n18450) );
  BUF_X1 U418 ( .A(n19076), .Z(n18447) );
  BUF_X1 U419 ( .A(n19074), .Z(n18444) );
  BUF_X1 U420 ( .A(n19120), .Z(n18513) );
  BUF_X1 U421 ( .A(n19118), .Z(n18510) );
  BUF_X1 U422 ( .A(n19116), .Z(n18507) );
  BUF_X1 U423 ( .A(n19114), .Z(n18504) );
  BUF_X1 U424 ( .A(n19112), .Z(n18501) );
  BUF_X1 U425 ( .A(n19110), .Z(n18498) );
  BUF_X1 U426 ( .A(n19108), .Z(n18495) );
  BUF_X1 U427 ( .A(n19106), .Z(n18492) );
  BUF_X1 U428 ( .A(n19072), .Z(n18441) );
  BUF_X1 U429 ( .A(n19070), .Z(n18438) );
  BUF_X1 U430 ( .A(n19068), .Z(n18435) );
  BUF_X1 U431 ( .A(n19066), .Z(n18432) );
  BUF_X1 U432 ( .A(n19064), .Z(n18429) );
  BUF_X1 U433 ( .A(n19062), .Z(n18426) );
  BUF_X1 U434 ( .A(n19060), .Z(n18423) );
  BUF_X1 U435 ( .A(n19058), .Z(n18420) );
  BUF_X1 U436 ( .A(n1631), .Z(n18545) );
  BUF_X1 U437 ( .A(n1641), .Z(n18521) );
  BUF_X1 U438 ( .A(n1631), .Z(n18546) );
  BUF_X1 U439 ( .A(n1641), .Z(n18522) );
  BUF_X1 U440 ( .A(n1006), .Z(n18654) );
  BUF_X1 U441 ( .A(n1011), .Z(n18642) );
  BUF_X1 U442 ( .A(n1016), .Z(n18630) );
  BUF_X1 U443 ( .A(n1021), .Z(n18618) );
  BUF_X1 U444 ( .A(n982), .Z(n18702) );
  BUF_X1 U445 ( .A(n987), .Z(n18690) );
  BUF_X1 U446 ( .A(n992), .Z(n18678) );
  BUF_X1 U447 ( .A(n997), .Z(n18666) );
  BUF_X1 U448 ( .A(n1011), .Z(n18641) );
  BUF_X1 U449 ( .A(n1016), .Z(n18629) );
  BUF_X1 U450 ( .A(n1021), .Z(n18617) );
  BUF_X1 U451 ( .A(n982), .Z(n18701) );
  BUF_X1 U452 ( .A(n992), .Z(n18677) );
  BUF_X1 U453 ( .A(n987), .Z(n18689) );
  BUF_X1 U454 ( .A(n997), .Z(n18665) );
  BUF_X1 U455 ( .A(n1602), .Z(n18605) );
  BUF_X1 U456 ( .A(n1607), .Z(n18593) );
  BUF_X1 U457 ( .A(n1612), .Z(n18581) );
  BUF_X1 U458 ( .A(n1617), .Z(n18569) );
  BUF_X1 U459 ( .A(n1626), .Z(n18557) );
  BUF_X1 U460 ( .A(n1636), .Z(n18533) );
  BUF_X1 U461 ( .A(n1602), .Z(n18606) );
  BUF_X1 U462 ( .A(n1607), .Z(n18594) );
  BUF_X1 U463 ( .A(n1612), .Z(n18582) );
  BUF_X1 U464 ( .A(n1617), .Z(n18570) );
  BUF_X1 U465 ( .A(n1626), .Z(n18558) );
  BUF_X1 U466 ( .A(n1636), .Z(n18534) );
  BUF_X1 U467 ( .A(n1008), .Z(n18651) );
  BUF_X1 U468 ( .A(n1013), .Z(n18639) );
  BUF_X1 U469 ( .A(n1018), .Z(n18627) );
  BUF_X1 U470 ( .A(n1023), .Z(n18615) );
  BUF_X1 U471 ( .A(n984), .Z(n18699) );
  BUF_X1 U472 ( .A(n989), .Z(n18687) );
  BUF_X1 U473 ( .A(n994), .Z(n18675) );
  BUF_X1 U474 ( .A(n999), .Z(n18663) );
  BUF_X1 U475 ( .A(n1008), .Z(n18650) );
  BUF_X1 U476 ( .A(n1013), .Z(n18638) );
  BUF_X1 U477 ( .A(n1018), .Z(n18626) );
  BUF_X1 U478 ( .A(n1023), .Z(n18614) );
  BUF_X1 U479 ( .A(n984), .Z(n18698) );
  BUF_X1 U480 ( .A(n994), .Z(n18674) );
  BUF_X1 U481 ( .A(n989), .Z(n18686) );
  BUF_X1 U482 ( .A(n999), .Z(n18662) );
  BUF_X1 U483 ( .A(n1604), .Z(n18602) );
  BUF_X1 U484 ( .A(n1609), .Z(n18590) );
  BUF_X1 U485 ( .A(n1614), .Z(n18578) );
  BUF_X1 U486 ( .A(n1619), .Z(n18566) );
  BUF_X1 U487 ( .A(n1628), .Z(n18554) );
  BUF_X1 U488 ( .A(n1638), .Z(n18530) );
  BUF_X1 U489 ( .A(n1633), .Z(n18542) );
  BUF_X1 U490 ( .A(n1643), .Z(n18518) );
  BUF_X1 U491 ( .A(n1604), .Z(n18603) );
  BUF_X1 U492 ( .A(n1609), .Z(n18591) );
  BUF_X1 U493 ( .A(n1614), .Z(n18579) );
  BUF_X1 U494 ( .A(n1619), .Z(n18567) );
  BUF_X1 U495 ( .A(n1628), .Z(n18555) );
  BUF_X1 U496 ( .A(n1638), .Z(n18531) );
  BUF_X1 U497 ( .A(n1633), .Z(n18543) );
  BUF_X1 U498 ( .A(n1643), .Z(n18519) );
  BUF_X1 U499 ( .A(n1630), .Z(n18548) );
  BUF_X1 U500 ( .A(n1640), .Z(n18524) );
  BUF_X1 U501 ( .A(n1630), .Z(n18549) );
  BUF_X1 U502 ( .A(n1640), .Z(n18525) );
  BUF_X1 U503 ( .A(n1005), .Z(n18657) );
  BUF_X1 U504 ( .A(n1010), .Z(n18645) );
  BUF_X1 U505 ( .A(n1015), .Z(n18633) );
  BUF_X1 U506 ( .A(n1020), .Z(n18621) );
  BUF_X1 U507 ( .A(n981), .Z(n18705) );
  BUF_X1 U508 ( .A(n986), .Z(n18693) );
  BUF_X1 U509 ( .A(n991), .Z(n18681) );
  BUF_X1 U510 ( .A(n996), .Z(n18669) );
  BUF_X1 U511 ( .A(n1010), .Z(n18644) );
  BUF_X1 U512 ( .A(n1015), .Z(n18632) );
  BUF_X1 U513 ( .A(n1020), .Z(n18620) );
  BUF_X1 U514 ( .A(n981), .Z(n18704) );
  BUF_X1 U515 ( .A(n991), .Z(n18680) );
  BUF_X1 U516 ( .A(n986), .Z(n18692) );
  BUF_X1 U517 ( .A(n996), .Z(n18668) );
  BUF_X1 U518 ( .A(n1601), .Z(n18608) );
  BUF_X1 U519 ( .A(n1606), .Z(n18596) );
  BUF_X1 U520 ( .A(n1611), .Z(n18584) );
  BUF_X1 U521 ( .A(n1616), .Z(n18572) );
  BUF_X1 U522 ( .A(n1625), .Z(n18560) );
  BUF_X1 U523 ( .A(n1635), .Z(n18536) );
  BUF_X1 U524 ( .A(n1601), .Z(n18609) );
  BUF_X1 U525 ( .A(n1606), .Z(n18597) );
  BUF_X1 U526 ( .A(n1611), .Z(n18585) );
  BUF_X1 U527 ( .A(n1616), .Z(n18573) );
  BUF_X1 U528 ( .A(n1625), .Z(n18561) );
  BUF_X1 U529 ( .A(n1635), .Z(n18537) );
  BUF_X1 U530 ( .A(n1006), .Z(n18653) );
  BUF_X1 U531 ( .A(n1005), .Z(n18656) );
  BUF_X1 U532 ( .A(n1009), .Z(n18648) );
  BUF_X1 U533 ( .A(n1014), .Z(n18636) );
  BUF_X1 U534 ( .A(n1019), .Z(n18624) );
  BUF_X1 U535 ( .A(n1024), .Z(n18612) );
  BUF_X1 U536 ( .A(n985), .Z(n18696) );
  BUF_X1 U537 ( .A(n990), .Z(n18684) );
  BUF_X1 U538 ( .A(n995), .Z(n18672) );
  BUF_X1 U539 ( .A(n1000), .Z(n18660) );
  BUF_X1 U540 ( .A(n1009), .Z(n18647) );
  BUF_X1 U541 ( .A(n1014), .Z(n18635) );
  BUF_X1 U542 ( .A(n1019), .Z(n18623) );
  BUF_X1 U543 ( .A(n1024), .Z(n18611) );
  BUF_X1 U544 ( .A(n985), .Z(n18695) );
  BUF_X1 U545 ( .A(n990), .Z(n18683) );
  BUF_X1 U546 ( .A(n995), .Z(n18671) );
  BUF_X1 U547 ( .A(n1000), .Z(n18659) );
  BUF_X1 U548 ( .A(n1605), .Z(n18600) );
  BUF_X1 U549 ( .A(n1610), .Z(n18588) );
  BUF_X1 U550 ( .A(n1615), .Z(n18576) );
  BUF_X1 U551 ( .A(n1620), .Z(n18564) );
  BUF_X1 U552 ( .A(n1629), .Z(n18552) );
  BUF_X1 U553 ( .A(n1639), .Z(n18528) );
  BUF_X1 U554 ( .A(n1634), .Z(n18540) );
  BUF_X1 U555 ( .A(n1644), .Z(n18516) );
  BUF_X1 U556 ( .A(n1605), .Z(n18599) );
  BUF_X1 U557 ( .A(n1610), .Z(n18587) );
  BUF_X1 U558 ( .A(n1615), .Z(n18575) );
  BUF_X1 U559 ( .A(n1620), .Z(n18563) );
  BUF_X1 U560 ( .A(n1629), .Z(n18551) );
  BUF_X1 U561 ( .A(n1639), .Z(n18527) );
  BUF_X1 U562 ( .A(n1634), .Z(n18539) );
  BUF_X1 U563 ( .A(n1644), .Z(n18515) );
  BUF_X1 U564 ( .A(n1631), .Z(n18547) );
  BUF_X1 U565 ( .A(n1641), .Z(n18523) );
  BUF_X1 U566 ( .A(n1006), .Z(n18655) );
  BUF_X1 U567 ( .A(n1011), .Z(n18643) );
  BUF_X1 U568 ( .A(n1016), .Z(n18631) );
  BUF_X1 U569 ( .A(n1021), .Z(n18619) );
  BUF_X1 U570 ( .A(n982), .Z(n18703) );
  BUF_X1 U571 ( .A(n987), .Z(n18691) );
  BUF_X1 U572 ( .A(n992), .Z(n18679) );
  BUF_X1 U573 ( .A(n997), .Z(n18667) );
  BUF_X1 U574 ( .A(n1607), .Z(n18595) );
  BUF_X1 U575 ( .A(n1602), .Z(n18607) );
  BUF_X1 U576 ( .A(n1612), .Z(n18583) );
  BUF_X1 U577 ( .A(n1617), .Z(n18571) );
  BUF_X1 U578 ( .A(n1626), .Z(n18559) );
  BUF_X1 U579 ( .A(n1636), .Z(n18535) );
  BUF_X1 U580 ( .A(n1008), .Z(n18652) );
  BUF_X1 U581 ( .A(n1013), .Z(n18640) );
  BUF_X1 U582 ( .A(n1023), .Z(n18616) );
  BUF_X1 U583 ( .A(n989), .Z(n18688) );
  BUF_X1 U584 ( .A(n1018), .Z(n18628) );
  BUF_X1 U585 ( .A(n984), .Z(n18700) );
  BUF_X1 U586 ( .A(n994), .Z(n18676) );
  BUF_X1 U587 ( .A(n999), .Z(n18664) );
  BUF_X1 U588 ( .A(n1604), .Z(n18604) );
  BUF_X1 U589 ( .A(n1609), .Z(n18592) );
  BUF_X1 U590 ( .A(n1614), .Z(n18580) );
  BUF_X1 U591 ( .A(n1619), .Z(n18568) );
  BUF_X1 U592 ( .A(n1628), .Z(n18556) );
  BUF_X1 U593 ( .A(n1638), .Z(n18532) );
  BUF_X1 U594 ( .A(n1633), .Z(n18544) );
  BUF_X1 U595 ( .A(n1643), .Z(n18520) );
  BUF_X1 U596 ( .A(n1630), .Z(n18550) );
  BUF_X1 U597 ( .A(n1640), .Z(n18526) );
  BUF_X1 U598 ( .A(n1005), .Z(n18658) );
  BUF_X1 U599 ( .A(n1606), .Z(n18598) );
  BUF_X1 U600 ( .A(n1010), .Z(n18646) );
  BUF_X1 U601 ( .A(n1015), .Z(n18634) );
  BUF_X1 U602 ( .A(n1020), .Z(n18622) );
  BUF_X1 U603 ( .A(n981), .Z(n18706) );
  BUF_X1 U604 ( .A(n986), .Z(n18694) );
  BUF_X1 U605 ( .A(n991), .Z(n18682) );
  BUF_X1 U606 ( .A(n996), .Z(n18670) );
  BUF_X1 U607 ( .A(n1601), .Z(n18610) );
  BUF_X1 U608 ( .A(n1611), .Z(n18586) );
  BUF_X1 U609 ( .A(n1616), .Z(n18574) );
  BUF_X1 U610 ( .A(n1625), .Z(n18562) );
  BUF_X1 U611 ( .A(n1635), .Z(n18538) );
  BUF_X1 U612 ( .A(n1014), .Z(n18637) );
  BUF_X1 U613 ( .A(n985), .Z(n18697) );
  BUF_X1 U614 ( .A(n990), .Z(n18685) );
  BUF_X1 U615 ( .A(n1009), .Z(n18649) );
  BUF_X1 U616 ( .A(n1019), .Z(n18625) );
  BUF_X1 U617 ( .A(n1024), .Z(n18613) );
  BUF_X1 U618 ( .A(n995), .Z(n18673) );
  BUF_X1 U619 ( .A(n1000), .Z(n18661) );
  BUF_X1 U620 ( .A(n1629), .Z(n18553) );
  BUF_X1 U621 ( .A(n1639), .Z(n18529) );
  BUF_X1 U622 ( .A(n1634), .Z(n18541) );
  BUF_X1 U623 ( .A(n1644), .Z(n18517) );
  BUF_X1 U624 ( .A(n1605), .Z(n18601) );
  BUF_X1 U625 ( .A(n1610), .Z(n18589) );
  BUF_X1 U626 ( .A(n1615), .Z(n18577) );
  BUF_X1 U627 ( .A(n1620), .Z(n18565) );
  BUF_X1 U628 ( .A(n898), .Z(n19053) );
  BUF_X1 U629 ( .A(n898), .Z(n19052) );
  BUF_X1 U630 ( .A(n898), .Z(n19051) );
  BUF_X1 U631 ( .A(n898), .Z(n19050) );
  BUF_X1 U632 ( .A(n898), .Z(n19049) );
  BUF_X1 U633 ( .A(n898), .Z(n19048) );
  BUF_X1 U634 ( .A(n19104), .Z(n18490) );
  BUF_X1 U635 ( .A(n19102), .Z(n18487) );
  BUF_X1 U636 ( .A(n19100), .Z(n18484) );
  BUF_X1 U637 ( .A(n19098), .Z(n18481) );
  BUF_X1 U638 ( .A(n19096), .Z(n18478) );
  BUF_X1 U639 ( .A(n19094), .Z(n18475) );
  BUF_X1 U640 ( .A(n19092), .Z(n18472) );
  BUF_X1 U641 ( .A(n19090), .Z(n18469) );
  BUF_X1 U642 ( .A(n19088), .Z(n18466) );
  BUF_X1 U643 ( .A(n19086), .Z(n18463) );
  BUF_X1 U644 ( .A(n19084), .Z(n18460) );
  BUF_X1 U645 ( .A(n19082), .Z(n18457) );
  BUF_X1 U646 ( .A(n19080), .Z(n18454) );
  BUF_X1 U647 ( .A(n19078), .Z(n18451) );
  BUF_X1 U648 ( .A(n19076), .Z(n18448) );
  BUF_X1 U649 ( .A(n19074), .Z(n18445) );
  BUF_X1 U650 ( .A(n19072), .Z(n18442) );
  BUF_X1 U651 ( .A(n19070), .Z(n18439) );
  BUF_X1 U652 ( .A(n19068), .Z(n18436) );
  BUF_X1 U653 ( .A(n19066), .Z(n18433) );
  BUF_X1 U654 ( .A(n19064), .Z(n18430) );
  BUF_X1 U655 ( .A(n19062), .Z(n18427) );
  BUF_X1 U656 ( .A(n19060), .Z(n18424) );
  BUF_X1 U657 ( .A(n19058), .Z(n18421) );
  BUF_X1 U658 ( .A(n19120), .Z(n18514) );
  BUF_X1 U659 ( .A(n19118), .Z(n18511) );
  BUF_X1 U660 ( .A(n19116), .Z(n18508) );
  BUF_X1 U661 ( .A(n19114), .Z(n18505) );
  BUF_X1 U662 ( .A(n19112), .Z(n18502) );
  BUF_X1 U663 ( .A(n19110), .Z(n18499) );
  BUF_X1 U664 ( .A(n19108), .Z(n18496) );
  BUF_X1 U665 ( .A(n19106), .Z(n18493) );
  BUF_X1 U666 ( .A(n904), .Z(n19030) );
  BUF_X1 U667 ( .A(n904), .Z(n19031) );
  BUF_X1 U668 ( .A(n904), .Z(n19032) );
  BUF_X1 U669 ( .A(n904), .Z(n19033) );
  BUF_X1 U670 ( .A(n904), .Z(n19028) );
  BUF_X1 U671 ( .A(n904), .Z(n19029) );
  BUF_X1 U672 ( .A(n898), .Z(n19054) );
  BUF_X1 U673 ( .A(n904), .Z(n19034) );
  INV_X1 U674 ( .A(n19055), .ZN(n19057) );
  NOR3_X1 U675 ( .A1(n19125), .A2(n19124), .A3(n19126), .ZN(n961) );
  NOR3_X1 U676 ( .A1(n19917), .A2(n19914), .A3(n19913), .ZN(n1575) );
  AND3_X1 U677 ( .A1(n19123), .A2(n19122), .A3(n970), .ZN(n943) );
  NAND2_X1 U678 ( .A1(n1576), .A2(n1583), .ZN(n1011) );
  NAND2_X1 U679 ( .A1(n1576), .A2(n1586), .ZN(n1020) );
  NAND2_X1 U680 ( .A1(n1576), .A2(n1574), .ZN(n982) );
  NAND2_X1 U681 ( .A1(n1579), .A2(n1574), .ZN(n996) );
  NAND2_X1 U682 ( .A1(n1577), .A2(n1586), .ZN(n1021) );
  NAND2_X1 U683 ( .A1(n1577), .A2(n1573), .ZN(n981) );
  NAND2_X1 U684 ( .A1(n1572), .A2(n1586), .ZN(n1015) );
  AOI22_X1 U685 ( .A1(n18662), .A2(n19888), .B1(n18661), .B2(n19542), .ZN(
        n1585) );
  AOI22_X1 U686 ( .A1(n18662), .A2(n19910), .B1(n18660), .B2(n19532), .ZN(
        n1394) );
  AOI22_X1 U687 ( .A1(n18662), .A2(n19909), .B1(n18660), .B2(n19531), .ZN(
        n1376) );
  AOI22_X1 U688 ( .A1(n18663), .A2(n19908), .B1(n18660), .B2(n19530), .ZN(
        n1358) );
  AOI22_X1 U689 ( .A1(n18663), .A2(n19903), .B1(n18660), .B2(n19525), .ZN(
        n1268) );
  AOI22_X1 U690 ( .A1(n18663), .A2(n19902), .B1(n18660), .B2(n19524), .ZN(
        n1250) );
  AOI22_X1 U691 ( .A1(n18663), .A2(n19901), .B1(n18660), .B2(n19523), .ZN(
        n1232) );
  AOI22_X1 U692 ( .A1(n18662), .A2(n19887), .B1(n18661), .B2(n19541), .ZN(
        n1556) );
  AOI22_X1 U693 ( .A1(n18663), .A2(n19907), .B1(n18660), .B2(n19529), .ZN(
        n1340) );
  AOI22_X1 U694 ( .A1(n18663), .A2(n19906), .B1(n18660), .B2(n19528), .ZN(
        n1322) );
  AOI22_X1 U695 ( .A1(n18663), .A2(n19905), .B1(n18660), .B2(n19527), .ZN(
        n1304) );
  AOI22_X1 U696 ( .A1(n18663), .A2(n19904), .B1(n18660), .B2(n19526), .ZN(
        n1286) );
  AOI22_X1 U697 ( .A1(n18663), .A2(n19900), .B1(n18659), .B2(n19522), .ZN(
        n1214) );
  AOI22_X1 U698 ( .A1(n18663), .A2(n19899), .B1(n18659), .B2(n19521), .ZN(
        n1196) );
  AOI22_X1 U699 ( .A1(n18663), .A2(n19898), .B1(n18659), .B2(n19520), .ZN(
        n1178) );
  AOI22_X1 U700 ( .A1(n18663), .A2(n19897), .B1(n18659), .B2(n19519), .ZN(
        n1160) );
  AOI22_X1 U701 ( .A1(n18662), .A2(n19882), .B1(n18661), .B2(n19536), .ZN(
        n1466) );
  AOI22_X1 U702 ( .A1(n18662), .A2(n19881), .B1(n18661), .B2(n19535), .ZN(
        n1448) );
  AOI22_X1 U703 ( .A1(n18662), .A2(n19912), .B1(n18660), .B2(n19534), .ZN(
        n1430) );
  AOI22_X1 U704 ( .A1(n18662), .A2(n19911), .B1(n18660), .B2(n19533), .ZN(
        n1412) );
  AOI22_X1 U705 ( .A1(n18662), .A2(n19885), .B1(n18661), .B2(n19539), .ZN(
        n1520) );
  AOI22_X1 U706 ( .A1(n18664), .A2(n19889), .B1(n18659), .B2(n19463), .ZN(n998) );
  AOI22_X1 U707 ( .A1(n18662), .A2(n19884), .B1(n18661), .B2(n19538), .ZN(
        n1502) );
  AOI22_X1 U708 ( .A1(n18662), .A2(n19883), .B1(n18661), .B2(n19537), .ZN(
        n1484) );
  AOI22_X1 U709 ( .A1(n18664), .A2(n19892), .B1(n18659), .B2(n19466), .ZN(
        n1070) );
  AOI22_X1 U710 ( .A1(n18664), .A2(n19891), .B1(n18659), .B2(n19465), .ZN(
        n1052) );
  AOI22_X1 U711 ( .A1(n18662), .A2(n19886), .B1(n18661), .B2(n19540), .ZN(
        n1538) );
  AOI22_X1 U712 ( .A1(n18664), .A2(n19890), .B1(n18659), .B2(n19464), .ZN(
        n1034) );
  AOI22_X1 U713 ( .A1(n18664), .A2(n19896), .B1(n18659), .B2(n19470), .ZN(
        n1142) );
  AOI22_X1 U714 ( .A1(n18664), .A2(n19895), .B1(n18659), .B2(n19469), .ZN(
        n1124) );
  AOI22_X1 U715 ( .A1(n18664), .A2(n19894), .B1(n18659), .B2(n19468), .ZN(
        n1106) );
  AOI22_X1 U716 ( .A1(n18664), .A2(n19893), .B1(n18659), .B2(n19467), .ZN(
        n1088) );
  OAI22_X1 U717 ( .A1(n18488), .A2(n18939), .B1(n18942), .B2(n19880), .ZN(
        n3826) );
  OAI22_X1 U718 ( .A1(n18485), .A2(n18939), .B1(n18942), .B2(n19879), .ZN(
        n3810) );
  OAI22_X1 U719 ( .A1(n18482), .A2(n18939), .B1(n18942), .B2(n19878), .ZN(
        n3794) );
  OAI22_X1 U720 ( .A1(n18479), .A2(n18939), .B1(n18942), .B2(n19877), .ZN(
        n3778) );
  OAI22_X1 U721 ( .A1(n18476), .A2(n18939), .B1(n18943), .B2(n19876), .ZN(
        n3762) );
  OAI22_X1 U722 ( .A1(n18473), .A2(n18939), .B1(n18943), .B2(n19875), .ZN(
        n3746) );
  OAI22_X1 U723 ( .A1(n18470), .A2(n18939), .B1(n18943), .B2(n19874), .ZN(
        n3730) );
  OAI22_X1 U724 ( .A1(n18467), .A2(n18939), .B1(n18943), .B2(n19873), .ZN(
        n3714) );
  OAI22_X1 U725 ( .A1(n18464), .A2(n18939), .B1(n18944), .B2(n19872), .ZN(
        n3698) );
  OAI22_X1 U726 ( .A1(n18461), .A2(n18939), .B1(n18944), .B2(n19871), .ZN(
        n3682) );
  OAI22_X1 U727 ( .A1(n18458), .A2(n18939), .B1(n18944), .B2(n19870), .ZN(
        n3666) );
  OAI22_X1 U728 ( .A1(n18455), .A2(n18939), .B1(n18944), .B2(n19869), .ZN(
        n3650) );
  OAI22_X1 U729 ( .A1(n18452), .A2(n18938), .B1(n18945), .B2(n19868), .ZN(
        n3634) );
  OAI22_X1 U730 ( .A1(n18449), .A2(n18938), .B1(n18945), .B2(n19867), .ZN(
        n3618) );
  OAI22_X1 U731 ( .A1(n18446), .A2(n18938), .B1(n18945), .B2(n19866), .ZN(
        n3602) );
  OAI22_X1 U732 ( .A1(n18443), .A2(n18938), .B1(n18945), .B2(n19865), .ZN(
        n3586) );
  OAI22_X1 U733 ( .A1(n18440), .A2(n18938), .B1(n18946), .B2(n19864), .ZN(
        n3570) );
  OAI22_X1 U734 ( .A1(n18437), .A2(n18938), .B1(n18946), .B2(n19863), .ZN(
        n3554) );
  OAI22_X1 U735 ( .A1(n18434), .A2(n18938), .B1(n18946), .B2(n19862), .ZN(
        n3538) );
  OAI22_X1 U736 ( .A1(n18431), .A2(n18938), .B1(n18946), .B2(n19861), .ZN(
        n3522) );
  OAI22_X1 U737 ( .A1(n18428), .A2(n18938), .B1(n18947), .B2(n19860), .ZN(
        n3506) );
  OAI22_X1 U738 ( .A1(n18425), .A2(n18938), .B1(n18947), .B2(n19859), .ZN(
        n3490) );
  OAI22_X1 U739 ( .A1(n18422), .A2(n18938), .B1(n18947), .B2(n19858), .ZN(
        n3474) );
  OAI22_X1 U740 ( .A1(n18419), .A2(n18938), .B1(n18947), .B2(n19857), .ZN(
        n3458) );
  OAI22_X1 U741 ( .A1(n18488), .A2(n18983), .B1(n18986), .B2(n19856), .ZN(
        n3830) );
  OAI22_X1 U742 ( .A1(n18485), .A2(n18983), .B1(n18986), .B2(n19855), .ZN(
        n3814) );
  OAI22_X1 U743 ( .A1(n18482), .A2(n18983), .B1(n18986), .B2(n19854), .ZN(
        n3798) );
  OAI22_X1 U744 ( .A1(n18479), .A2(n18983), .B1(n18986), .B2(n19853), .ZN(
        n3782) );
  OAI22_X1 U745 ( .A1(n18476), .A2(n18983), .B1(n18987), .B2(n19852), .ZN(
        n3766) );
  OAI22_X1 U746 ( .A1(n18473), .A2(n18983), .B1(n18987), .B2(n19851), .ZN(
        n3750) );
  OAI22_X1 U747 ( .A1(n18470), .A2(n18983), .B1(n18987), .B2(n19850), .ZN(
        n3734) );
  OAI22_X1 U748 ( .A1(n18467), .A2(n18983), .B1(n18987), .B2(n19849), .ZN(
        n3718) );
  OAI22_X1 U749 ( .A1(n18464), .A2(n18983), .B1(n18988), .B2(n19848), .ZN(
        n3702) );
  OAI22_X1 U750 ( .A1(n18461), .A2(n18983), .B1(n18988), .B2(n19847), .ZN(
        n3686) );
  OAI22_X1 U751 ( .A1(n18458), .A2(n18983), .B1(n18988), .B2(n19846), .ZN(
        n3670) );
  OAI22_X1 U752 ( .A1(n18455), .A2(n18983), .B1(n18988), .B2(n19845), .ZN(
        n3654) );
  OAI22_X1 U753 ( .A1(n18452), .A2(n18982), .B1(n18989), .B2(n19844), .ZN(
        n3638) );
  OAI22_X1 U754 ( .A1(n18449), .A2(n18982), .B1(n18989), .B2(n19843), .ZN(
        n3622) );
  OAI22_X1 U755 ( .A1(n18446), .A2(n18982), .B1(n18989), .B2(n19842), .ZN(
        n3606) );
  OAI22_X1 U756 ( .A1(n18443), .A2(n18982), .B1(n18989), .B2(n19841), .ZN(
        n3590) );
  OAI22_X1 U757 ( .A1(n18440), .A2(n18982), .B1(n18990), .B2(n19840), .ZN(
        n3574) );
  OAI22_X1 U758 ( .A1(n18437), .A2(n18982), .B1(n18990), .B2(n19839), .ZN(
        n3558) );
  OAI22_X1 U759 ( .A1(n18434), .A2(n18982), .B1(n18990), .B2(n19838), .ZN(
        n3542) );
  OAI22_X1 U760 ( .A1(n18431), .A2(n18982), .B1(n18990), .B2(n19837), .ZN(
        n3526) );
  OAI22_X1 U761 ( .A1(n18428), .A2(n18982), .B1(n18991), .B2(n19836), .ZN(
        n3510) );
  OAI22_X1 U762 ( .A1(n18425), .A2(n18982), .B1(n18991), .B2(n19835), .ZN(
        n3494) );
  OAI22_X1 U763 ( .A1(n18422), .A2(n18982), .B1(n18991), .B2(n19834), .ZN(
        n3478) );
  OAI22_X1 U764 ( .A1(n18419), .A2(n18982), .B1(n18991), .B2(n19833), .ZN(
        n3462) );
  OAI22_X1 U765 ( .A1(n18513), .A2(n18861), .B1(n18870), .B2(n19832), .ZN(
        n3358) );
  OAI22_X1 U766 ( .A1(n18510), .A2(n18861), .B1(n18870), .B2(n19831), .ZN(
        n3359) );
  OAI22_X1 U767 ( .A1(n18507), .A2(n18861), .B1(n18870), .B2(n19830), .ZN(
        n3360) );
  OAI22_X1 U768 ( .A1(n18504), .A2(n18861), .B1(n18870), .B2(n19829), .ZN(
        n3361) );
  OAI22_X1 U769 ( .A1(n18501), .A2(n18861), .B1(n18869), .B2(n19828), .ZN(
        n3362) );
  OAI22_X1 U770 ( .A1(n18498), .A2(n18861), .B1(n18869), .B2(n19827), .ZN(
        n3363) );
  OAI22_X1 U771 ( .A1(n18495), .A2(n18861), .B1(n18869), .B2(n19826), .ZN(
        n3364) );
  OAI22_X1 U772 ( .A1(n18492), .A2(n18861), .B1(n18869), .B2(n19825), .ZN(
        n3365) );
  OAI22_X1 U773 ( .A1(n18489), .A2(n18861), .B1(n18868), .B2(n19824), .ZN(
        n3366) );
  OAI22_X1 U774 ( .A1(n18486), .A2(n18861), .B1(n18868), .B2(n19823), .ZN(
        n3367) );
  OAI22_X1 U775 ( .A1(n18513), .A2(n18817), .B1(n18826), .B2(n19822), .ZN(
        n3230) );
  OAI22_X1 U776 ( .A1(n18510), .A2(n18817), .B1(n18826), .B2(n19821), .ZN(
        n3231) );
  OAI22_X1 U777 ( .A1(n18507), .A2(n18817), .B1(n18826), .B2(n19820), .ZN(
        n3232) );
  OAI22_X1 U778 ( .A1(n18504), .A2(n18817), .B1(n18826), .B2(n19819), .ZN(
        n3233) );
  OAI22_X1 U779 ( .A1(n18501), .A2(n18817), .B1(n18825), .B2(n19818), .ZN(
        n3234) );
  OAI22_X1 U780 ( .A1(n18498), .A2(n18817), .B1(n18825), .B2(n19817), .ZN(
        n3235) );
  OAI22_X1 U781 ( .A1(n18495), .A2(n18817), .B1(n18825), .B2(n19816), .ZN(
        n3236) );
  OAI22_X1 U782 ( .A1(n18492), .A2(n18817), .B1(n18825), .B2(n19815), .ZN(
        n3237) );
  OAI22_X1 U783 ( .A1(n18489), .A2(n18817), .B1(n18824), .B2(n19814), .ZN(
        n3238) );
  OAI22_X1 U784 ( .A1(n18486), .A2(n18817), .B1(n18824), .B2(n19813), .ZN(
        n3239) );
  OAI22_X1 U785 ( .A1(n18483), .A2(n18817), .B1(n18824), .B2(n19812), .ZN(
        n3240) );
  OAI22_X1 U786 ( .A1(n18480), .A2(n18817), .B1(n18824), .B2(n19811), .ZN(
        n3241) );
  OAI22_X1 U787 ( .A1(n18477), .A2(n18818), .B1(n18823), .B2(n19810), .ZN(
        n3242) );
  OAI22_X1 U788 ( .A1(n18474), .A2(n18818), .B1(n18823), .B2(n19809), .ZN(
        n3243) );
  OAI22_X1 U789 ( .A1(n18471), .A2(n18818), .B1(n18823), .B2(n19808), .ZN(
        n3244) );
  OAI22_X1 U790 ( .A1(n18468), .A2(n18818), .B1(n18823), .B2(n19807), .ZN(
        n3245) );
  OAI22_X1 U791 ( .A1(n18465), .A2(n18818), .B1(n18822), .B2(n19806), .ZN(
        n3246) );
  OAI22_X1 U792 ( .A1(n18462), .A2(n18818), .B1(n18822), .B2(n19805), .ZN(
        n3247) );
  OAI22_X1 U793 ( .A1(n18459), .A2(n18818), .B1(n18822), .B2(n19804), .ZN(
        n3248) );
  OAI22_X1 U794 ( .A1(n18456), .A2(n18818), .B1(n18822), .B2(n19803), .ZN(
        n3249) );
  OAI22_X1 U795 ( .A1(n18453), .A2(n18818), .B1(n18821), .B2(n19802), .ZN(
        n3250) );
  OAI22_X1 U796 ( .A1(n18450), .A2(n18818), .B1(n18821), .B2(n19801), .ZN(
        n3251) );
  OAI22_X1 U797 ( .A1(n18447), .A2(n18818), .B1(n18821), .B2(n19800), .ZN(
        n3252) );
  OAI22_X1 U798 ( .A1(n18444), .A2(n18818), .B1(n18821), .B2(n19799), .ZN(
        n3253) );
  OAI22_X1 U799 ( .A1(n18513), .A2(n18773), .B1(n18782), .B2(n19774), .ZN(
        n3102) );
  OAI22_X1 U800 ( .A1(n18510), .A2(n18773), .B1(n18782), .B2(n19773), .ZN(
        n3103) );
  OAI22_X1 U801 ( .A1(n18507), .A2(n18773), .B1(n18782), .B2(n19772), .ZN(
        n3104) );
  OAI22_X1 U802 ( .A1(n18504), .A2(n18773), .B1(n18782), .B2(n19771), .ZN(
        n3105) );
  OAI22_X1 U803 ( .A1(n18501), .A2(n18773), .B1(n18781), .B2(n19770), .ZN(
        n3106) );
  OAI22_X1 U804 ( .A1(n18498), .A2(n18773), .B1(n18781), .B2(n19769), .ZN(
        n3107) );
  OAI22_X1 U805 ( .A1(n18495), .A2(n18773), .B1(n18781), .B2(n19768), .ZN(
        n3108) );
  OAI22_X1 U806 ( .A1(n18492), .A2(n18773), .B1(n18781), .B2(n19767), .ZN(
        n3109) );
  OAI22_X1 U807 ( .A1(n18489), .A2(n18773), .B1(n18780), .B2(n19766), .ZN(
        n3110) );
  OAI22_X1 U808 ( .A1(n18486), .A2(n18773), .B1(n18780), .B2(n19765), .ZN(
        n3111) );
  OAI22_X1 U809 ( .A1(n18483), .A2(n18773), .B1(n18780), .B2(n19764), .ZN(
        n3112) );
  OAI22_X1 U810 ( .A1(n18480), .A2(n18773), .B1(n18780), .B2(n19763), .ZN(
        n3113) );
  OAI22_X1 U811 ( .A1(n18477), .A2(n18774), .B1(n18779), .B2(n19762), .ZN(
        n3114) );
  OAI22_X1 U812 ( .A1(n18474), .A2(n18774), .B1(n18779), .B2(n19761), .ZN(
        n3115) );
  OAI22_X1 U813 ( .A1(n18471), .A2(n18774), .B1(n18779), .B2(n19760), .ZN(
        n3116) );
  OAI22_X1 U814 ( .A1(n18468), .A2(n18774), .B1(n18779), .B2(n19759), .ZN(
        n3117) );
  OAI22_X1 U815 ( .A1(n18465), .A2(n18774), .B1(n18778), .B2(n19758), .ZN(
        n3118) );
  OAI22_X1 U816 ( .A1(n18462), .A2(n18774), .B1(n18778), .B2(n19757), .ZN(
        n3119) );
  OAI22_X1 U817 ( .A1(n18459), .A2(n18774), .B1(n18778), .B2(n19756), .ZN(
        n3120) );
  OAI22_X1 U818 ( .A1(n18456), .A2(n18774), .B1(n18778), .B2(n19755), .ZN(
        n3121) );
  OAI22_X1 U819 ( .A1(n18453), .A2(n18774), .B1(n18777), .B2(n19754), .ZN(
        n3122) );
  OAI22_X1 U820 ( .A1(n18450), .A2(n18774), .B1(n18777), .B2(n19753), .ZN(
        n3123) );
  OAI22_X1 U821 ( .A1(n18447), .A2(n18774), .B1(n18777), .B2(n19752), .ZN(
        n3124) );
  OAI22_X1 U822 ( .A1(n18444), .A2(n18774), .B1(n18777), .B2(n19751), .ZN(
        n3125) );
  OAI22_X1 U823 ( .A1(n18488), .A2(n18961), .B1(n18964), .B2(n19750), .ZN(
        n3828) );
  OAI22_X1 U824 ( .A1(n18485), .A2(n18961), .B1(n18964), .B2(n19749), .ZN(
        n3812) );
  OAI22_X1 U825 ( .A1(n18482), .A2(n18961), .B1(n18964), .B2(n19748), .ZN(
        n3796) );
  OAI22_X1 U826 ( .A1(n18479), .A2(n18961), .B1(n18964), .B2(n19747), .ZN(
        n3780) );
  OAI22_X1 U827 ( .A1(n18476), .A2(n18961), .B1(n18965), .B2(n19746), .ZN(
        n3764) );
  OAI22_X1 U828 ( .A1(n18473), .A2(n18961), .B1(n18965), .B2(n19745), .ZN(
        n3748) );
  OAI22_X1 U829 ( .A1(n18470), .A2(n18961), .B1(n18965), .B2(n19744), .ZN(
        n3732) );
  OAI22_X1 U830 ( .A1(n18467), .A2(n18961), .B1(n18965), .B2(n19743), .ZN(
        n3716) );
  OAI22_X1 U831 ( .A1(n18464), .A2(n18961), .B1(n18966), .B2(n19742), .ZN(
        n3700) );
  OAI22_X1 U832 ( .A1(n18461), .A2(n18961), .B1(n18966), .B2(n19741), .ZN(
        n3684) );
  OAI22_X1 U833 ( .A1(n18458), .A2(n18961), .B1(n18966), .B2(n19740), .ZN(
        n3668) );
  OAI22_X1 U834 ( .A1(n18455), .A2(n18961), .B1(n18966), .B2(n19739), .ZN(
        n3652) );
  OAI22_X1 U835 ( .A1(n18452), .A2(n18960), .B1(n18967), .B2(n19738), .ZN(
        n3636) );
  OAI22_X1 U836 ( .A1(n18449), .A2(n18960), .B1(n18967), .B2(n19737), .ZN(
        n3620) );
  OAI22_X1 U837 ( .A1(n18446), .A2(n18960), .B1(n18967), .B2(n19736), .ZN(
        n3604) );
  OAI22_X1 U838 ( .A1(n18443), .A2(n18960), .B1(n18967), .B2(n19735), .ZN(
        n3588) );
  OAI22_X1 U839 ( .A1(n18440), .A2(n18960), .B1(n18968), .B2(n19734), .ZN(
        n3572) );
  OAI22_X1 U840 ( .A1(n18437), .A2(n18960), .B1(n18968), .B2(n19733), .ZN(
        n3556) );
  OAI22_X1 U841 ( .A1(n18434), .A2(n18960), .B1(n18968), .B2(n19732), .ZN(
        n3540) );
  OAI22_X1 U842 ( .A1(n18431), .A2(n18960), .B1(n18968), .B2(n19731), .ZN(
        n3524) );
  OAI22_X1 U843 ( .A1(n18428), .A2(n18960), .B1(n18969), .B2(n19730), .ZN(
        n3508) );
  OAI22_X1 U844 ( .A1(n18425), .A2(n18960), .B1(n18969), .B2(n19729), .ZN(
        n3492) );
  OAI22_X1 U845 ( .A1(n18422), .A2(n18960), .B1(n18969), .B2(n19728), .ZN(
        n3476) );
  OAI22_X1 U846 ( .A1(n18419), .A2(n18960), .B1(n18969), .B2(n19727), .ZN(
        n3460) );
  OAI22_X1 U847 ( .A1(n18513), .A2(n18828), .B1(n18837), .B2(n19726), .ZN(
        n3262) );
  OAI22_X1 U848 ( .A1(n18510), .A2(n18828), .B1(n18837), .B2(n19725), .ZN(
        n3263) );
  OAI22_X1 U849 ( .A1(n18507), .A2(n18828), .B1(n18837), .B2(n19724), .ZN(
        n3264) );
  OAI22_X1 U850 ( .A1(n18504), .A2(n18828), .B1(n18837), .B2(n19723), .ZN(
        n3265) );
  OAI22_X1 U851 ( .A1(n18501), .A2(n18828), .B1(n18836), .B2(n19722), .ZN(
        n3266) );
  OAI22_X1 U852 ( .A1(n18498), .A2(n18828), .B1(n18836), .B2(n19721), .ZN(
        n3267) );
  OAI22_X1 U853 ( .A1(n18495), .A2(n18828), .B1(n18836), .B2(n19720), .ZN(
        n3268) );
  OAI22_X1 U854 ( .A1(n18492), .A2(n18828), .B1(n18836), .B2(n19719), .ZN(
        n3269) );
  OAI22_X1 U855 ( .A1(n18489), .A2(n18828), .B1(n18835), .B2(n19718), .ZN(
        n3270) );
  OAI22_X1 U856 ( .A1(n18486), .A2(n18828), .B1(n18835), .B2(n19717), .ZN(
        n3271) );
  OAI22_X1 U857 ( .A1(n18483), .A2(n18828), .B1(n18835), .B2(n19716), .ZN(
        n3272) );
  OAI22_X1 U858 ( .A1(n18480), .A2(n18828), .B1(n18835), .B2(n19715), .ZN(
        n3273) );
  OAI22_X1 U859 ( .A1(n18477), .A2(n18829), .B1(n18834), .B2(n19714), .ZN(
        n3274) );
  OAI22_X1 U860 ( .A1(n18474), .A2(n18829), .B1(n18834), .B2(n19713), .ZN(
        n3275) );
  OAI22_X1 U861 ( .A1(n18471), .A2(n18829), .B1(n18834), .B2(n19712), .ZN(
        n3276) );
  OAI22_X1 U862 ( .A1(n18468), .A2(n18829), .B1(n18834), .B2(n19711), .ZN(
        n3277) );
  OAI22_X1 U863 ( .A1(n18465), .A2(n18829), .B1(n18833), .B2(n19710), .ZN(
        n3278) );
  OAI22_X1 U864 ( .A1(n18462), .A2(n18829), .B1(n18833), .B2(n19709), .ZN(
        n3279) );
  OAI22_X1 U865 ( .A1(n18459), .A2(n18829), .B1(n18833), .B2(n19708), .ZN(
        n3280) );
  OAI22_X1 U866 ( .A1(n18456), .A2(n18829), .B1(n18833), .B2(n19707), .ZN(
        n3281) );
  OAI22_X1 U867 ( .A1(n18453), .A2(n18829), .B1(n18832), .B2(n19706), .ZN(
        n3282) );
  OAI22_X1 U868 ( .A1(n18450), .A2(n18829), .B1(n18832), .B2(n19705), .ZN(
        n3283) );
  OAI22_X1 U869 ( .A1(n18447), .A2(n18829), .B1(n18832), .B2(n19704), .ZN(
        n3284) );
  OAI22_X1 U870 ( .A1(n18444), .A2(n18829), .B1(n18832), .B2(n19703), .ZN(
        n3285) );
  OAI22_X1 U871 ( .A1(n18512), .A2(n18939), .B1(n18940), .B2(n19678), .ZN(
        n3954) );
  OAI22_X1 U872 ( .A1(n18509), .A2(n18938), .B1(n18940), .B2(n19677), .ZN(
        n3938) );
  OAI22_X1 U873 ( .A1(n18506), .A2(n18939), .B1(n18940), .B2(n19676), .ZN(
        n3922) );
  OAI22_X1 U874 ( .A1(n18503), .A2(n18938), .B1(n18940), .B2(n19675), .ZN(
        n3906) );
  OAI22_X1 U875 ( .A1(n18500), .A2(n18939), .B1(n18941), .B2(n19674), .ZN(
        n3890) );
  OAI22_X1 U876 ( .A1(n18497), .A2(n18938), .B1(n18941), .B2(n19673), .ZN(
        n3874) );
  OAI22_X1 U877 ( .A1(n18494), .A2(n18939), .B1(n18941), .B2(n19672), .ZN(
        n3858) );
  OAI22_X1 U878 ( .A1(n18491), .A2(n18938), .B1(n18941), .B2(n19671), .ZN(
        n3842) );
  OAI22_X1 U879 ( .A1(n18512), .A2(n18983), .B1(n18984), .B2(n19670), .ZN(
        n3958) );
  OAI22_X1 U880 ( .A1(n18509), .A2(n18982), .B1(n18984), .B2(n19669), .ZN(
        n3942) );
  OAI22_X1 U881 ( .A1(n18506), .A2(n18983), .B1(n18984), .B2(n19668), .ZN(
        n3926) );
  OAI22_X1 U882 ( .A1(n18503), .A2(n18982), .B1(n18984), .B2(n19667), .ZN(
        n3910) );
  OAI22_X1 U883 ( .A1(n18500), .A2(n18983), .B1(n18985), .B2(n19666), .ZN(
        n3894) );
  OAI22_X1 U884 ( .A1(n18497), .A2(n18982), .B1(n18985), .B2(n19665), .ZN(
        n3878) );
  OAI22_X1 U885 ( .A1(n18494), .A2(n18983), .B1(n18985), .B2(n19664), .ZN(
        n3862) );
  OAI22_X1 U886 ( .A1(n18491), .A2(n18982), .B1(n18985), .B2(n19663), .ZN(
        n3846) );
  OAI22_X1 U887 ( .A1(n18441), .A2(n18861), .B1(n18867), .B2(n19662), .ZN(
        n3382) );
  OAI22_X1 U888 ( .A1(n18438), .A2(n18862), .B1(n18867), .B2(n19661), .ZN(
        n3383) );
  OAI22_X1 U889 ( .A1(n18435), .A2(n18861), .B1(n18867), .B2(n19660), .ZN(
        n3384) );
  OAI22_X1 U890 ( .A1(n18432), .A2(n18861), .B1(n18866), .B2(n19659), .ZN(
        n3385) );
  OAI22_X1 U891 ( .A1(n18429), .A2(n18862), .B1(n18868), .B2(n19658), .ZN(
        n3386) );
  OAI22_X1 U892 ( .A1(n18426), .A2(n18862), .B1(n18866), .B2(n19657), .ZN(
        n3387) );
  OAI22_X1 U893 ( .A1(n18423), .A2(n18861), .B1(n18867), .B2(n19656), .ZN(
        n3388) );
  OAI22_X1 U894 ( .A1(n18420), .A2(n18862), .B1(n18868), .B2(n19655), .ZN(
        n3389) );
  OAI22_X1 U895 ( .A1(n18441), .A2(n18817), .B1(n18820), .B2(n19654), .ZN(
        n3254) );
  OAI22_X1 U896 ( .A1(n18438), .A2(n18818), .B1(n18820), .B2(n19653), .ZN(
        n3255) );
  OAI22_X1 U897 ( .A1(n18435), .A2(n18817), .B1(n18820), .B2(n19652), .ZN(
        n3256) );
  OAI22_X1 U898 ( .A1(n18432), .A2(n18818), .B1(n18820), .B2(n19651), .ZN(
        n3257) );
  OAI22_X1 U899 ( .A1(n18429), .A2(n18817), .B1(n18819), .B2(n19650), .ZN(
        n3258) );
  OAI22_X1 U900 ( .A1(n18426), .A2(n18818), .B1(n18819), .B2(n19649), .ZN(
        n3259) );
  OAI22_X1 U901 ( .A1(n18423), .A2(n18817), .B1(n18819), .B2(n19648), .ZN(
        n3260) );
  OAI22_X1 U902 ( .A1(n18420), .A2(n18818), .B1(n18819), .B2(n19647), .ZN(
        n3261) );
  OAI22_X1 U903 ( .A1(n18441), .A2(n18773), .B1(n18776), .B2(n19638), .ZN(
        n3126) );
  OAI22_X1 U904 ( .A1(n18438), .A2(n18774), .B1(n18776), .B2(n19637), .ZN(
        n3127) );
  OAI22_X1 U905 ( .A1(n18435), .A2(n18773), .B1(n18776), .B2(n19636), .ZN(
        n3128) );
  OAI22_X1 U906 ( .A1(n18432), .A2(n18774), .B1(n18776), .B2(n19635), .ZN(
        n3129) );
  OAI22_X1 U907 ( .A1(n18429), .A2(n18773), .B1(n18775), .B2(n19634), .ZN(
        n3130) );
  OAI22_X1 U908 ( .A1(n18426), .A2(n18774), .B1(n18775), .B2(n19633), .ZN(
        n3131) );
  OAI22_X1 U909 ( .A1(n18423), .A2(n18773), .B1(n18775), .B2(n19632), .ZN(
        n3132) );
  OAI22_X1 U910 ( .A1(n18420), .A2(n18774), .B1(n18775), .B2(n19631), .ZN(
        n3133) );
  OAI22_X1 U911 ( .A1(n18512), .A2(n18961), .B1(n18962), .B2(n19630), .ZN(
        n3956) );
  OAI22_X1 U912 ( .A1(n18509), .A2(n18960), .B1(n18962), .B2(n19629), .ZN(
        n3940) );
  OAI22_X1 U913 ( .A1(n18506), .A2(n18961), .B1(n18962), .B2(n19628), .ZN(
        n3924) );
  OAI22_X1 U914 ( .A1(n18503), .A2(n18960), .B1(n18962), .B2(n19627), .ZN(
        n3908) );
  OAI22_X1 U915 ( .A1(n18500), .A2(n18961), .B1(n18963), .B2(n19626), .ZN(
        n3892) );
  OAI22_X1 U916 ( .A1(n18497), .A2(n18960), .B1(n18963), .B2(n19625), .ZN(
        n3876) );
  OAI22_X1 U917 ( .A1(n18494), .A2(n18961), .B1(n18963), .B2(n19624), .ZN(
        n3860) );
  OAI22_X1 U918 ( .A1(n18491), .A2(n18960), .B1(n18963), .B2(n19623), .ZN(
        n3844) );
  OAI22_X1 U919 ( .A1(n18441), .A2(n18828), .B1(n18831), .B2(n19622), .ZN(
        n3286) );
  OAI22_X1 U920 ( .A1(n18438), .A2(n18829), .B1(n18831), .B2(n19621), .ZN(
        n3287) );
  OAI22_X1 U921 ( .A1(n18435), .A2(n18828), .B1(n18831), .B2(n19620), .ZN(
        n3288) );
  OAI22_X1 U922 ( .A1(n18432), .A2(n18829), .B1(n18831), .B2(n19619), .ZN(
        n3289) );
  OAI22_X1 U923 ( .A1(n18429), .A2(n18828), .B1(n18830), .B2(n19618), .ZN(
        n3290) );
  OAI22_X1 U924 ( .A1(n18426), .A2(n18829), .B1(n18830), .B2(n19617), .ZN(
        n3291) );
  OAI22_X1 U925 ( .A1(n18423), .A2(n18828), .B1(n18830), .B2(n19616), .ZN(
        n3292) );
  OAI22_X1 U926 ( .A1(n18420), .A2(n18829), .B1(n18830), .B2(n19615), .ZN(
        n3293) );
  OAI22_X1 U927 ( .A1(n18512), .A2(n19004), .B1(n19013), .B2(n19606), .ZN(
        n9014) );
  OAI22_X1 U928 ( .A1(n18509), .A2(n19004), .B1(n19013), .B2(n19605), .ZN(
        n9015) );
  OAI22_X1 U929 ( .A1(n18506), .A2(n19004), .B1(n19013), .B2(n19604), .ZN(
        n9016) );
  OAI22_X1 U930 ( .A1(n18503), .A2(n19004), .B1(n19013), .B2(n19603), .ZN(
        n9017) );
  OAI22_X1 U931 ( .A1(n18500), .A2(n19004), .B1(n19012), .B2(n19602), .ZN(
        n9018) );
  OAI22_X1 U932 ( .A1(n18497), .A2(n19004), .B1(n19012), .B2(n19601), .ZN(
        n9019) );
  OAI22_X1 U933 ( .A1(n18494), .A2(n19004), .B1(n19012), .B2(n19600), .ZN(
        n9020) );
  OAI22_X1 U934 ( .A1(n18491), .A2(n19004), .B1(n19012), .B2(n19599), .ZN(
        n9021) );
  OAI22_X1 U935 ( .A1(n18488), .A2(n19004), .B1(n19011), .B2(n19598), .ZN(
        n9022) );
  OAI22_X1 U936 ( .A1(n18485), .A2(n19004), .B1(n19011), .B2(n19597), .ZN(
        n9023) );
  OAI22_X1 U937 ( .A1(n18482), .A2(n19004), .B1(n19011), .B2(n19596), .ZN(
        n9024) );
  OAI22_X1 U938 ( .A1(n18479), .A2(n19004), .B1(n19011), .B2(n19595), .ZN(
        n9025) );
  OAI22_X1 U939 ( .A1(n18476), .A2(n19005), .B1(n19010), .B2(n19594), .ZN(
        n9026) );
  OAI22_X1 U940 ( .A1(n18473), .A2(n19005), .B1(n19010), .B2(n19593), .ZN(
        n9027) );
  OAI22_X1 U941 ( .A1(n18470), .A2(n19005), .B1(n19010), .B2(n19592), .ZN(
        n9028) );
  OAI22_X1 U942 ( .A1(n18467), .A2(n19005), .B1(n19010), .B2(n19591), .ZN(
        n9029) );
  OAI22_X1 U943 ( .A1(n18464), .A2(n19005), .B1(n19009), .B2(n19590), .ZN(
        n9030) );
  OAI22_X1 U944 ( .A1(n18461), .A2(n19005), .B1(n19009), .B2(n19589), .ZN(
        n9031) );
  OAI22_X1 U945 ( .A1(n18458), .A2(n19005), .B1(n19009), .B2(n19588), .ZN(
        n9032) );
  OAI22_X1 U946 ( .A1(n18455), .A2(n19005), .B1(n19009), .B2(n19587), .ZN(
        n9033) );
  OAI22_X1 U947 ( .A1(n18452), .A2(n19005), .B1(n19008), .B2(n19586), .ZN(
        n9034) );
  OAI22_X1 U948 ( .A1(n18449), .A2(n19005), .B1(n19008), .B2(n19585), .ZN(
        n9035) );
  OAI22_X1 U949 ( .A1(n18446), .A2(n19005), .B1(n19008), .B2(n19584), .ZN(
        n9036) );
  OAI22_X1 U950 ( .A1(n18443), .A2(n19005), .B1(n19008), .B2(n19583), .ZN(
        n9037) );
  OAI22_X1 U951 ( .A1(n18488), .A2(n18950), .B1(n18953), .B2(n19582), .ZN(
        n3827) );
  OAI22_X1 U952 ( .A1(n18485), .A2(n18950), .B1(n18953), .B2(n19581), .ZN(
        n3811) );
  OAI22_X1 U953 ( .A1(n18482), .A2(n18950), .B1(n18953), .B2(n19580), .ZN(
        n3795) );
  OAI22_X1 U954 ( .A1(n18479), .A2(n18950), .B1(n18953), .B2(n19579), .ZN(
        n3779) );
  OAI22_X1 U955 ( .A1(n18476), .A2(n18950), .B1(n18954), .B2(n19578), .ZN(
        n3763) );
  OAI22_X1 U956 ( .A1(n18473), .A2(n18950), .B1(n18954), .B2(n19577), .ZN(
        n3747) );
  OAI22_X1 U957 ( .A1(n18470), .A2(n18950), .B1(n18954), .B2(n19576), .ZN(
        n3731) );
  OAI22_X1 U958 ( .A1(n18467), .A2(n18950), .B1(n18954), .B2(n19575), .ZN(
        n3715) );
  OAI22_X1 U959 ( .A1(n18464), .A2(n18950), .B1(n18955), .B2(n19574), .ZN(
        n3699) );
  OAI22_X1 U960 ( .A1(n18461), .A2(n18950), .B1(n18955), .B2(n19573), .ZN(
        n3683) );
  OAI22_X1 U961 ( .A1(n18458), .A2(n18950), .B1(n18955), .B2(n19572), .ZN(
        n3667) );
  OAI22_X1 U962 ( .A1(n18455), .A2(n18950), .B1(n18955), .B2(n19571), .ZN(
        n3651) );
  OAI22_X1 U963 ( .A1(n18452), .A2(n18949), .B1(n18956), .B2(n19570), .ZN(
        n3635) );
  OAI22_X1 U964 ( .A1(n18449), .A2(n18949), .B1(n18956), .B2(n19569), .ZN(
        n3619) );
  OAI22_X1 U965 ( .A1(n18446), .A2(n18949), .B1(n18956), .B2(n19568), .ZN(
        n3603) );
  OAI22_X1 U966 ( .A1(n18443), .A2(n18949), .B1(n18956), .B2(n19567), .ZN(
        n3587) );
  OAI22_X1 U967 ( .A1(n18440), .A2(n18949), .B1(n18957), .B2(n19566), .ZN(
        n3571) );
  OAI22_X1 U968 ( .A1(n18437), .A2(n18949), .B1(n18957), .B2(n19565), .ZN(
        n3555) );
  OAI22_X1 U969 ( .A1(n18434), .A2(n18949), .B1(n18957), .B2(n19564), .ZN(
        n3539) );
  OAI22_X1 U970 ( .A1(n18431), .A2(n18949), .B1(n18957), .B2(n19563), .ZN(
        n3523) );
  OAI22_X1 U971 ( .A1(n18428), .A2(n18949), .B1(n18958), .B2(n19562), .ZN(
        n3507) );
  OAI22_X1 U972 ( .A1(n18425), .A2(n18949), .B1(n18958), .B2(n19561), .ZN(
        n3491) );
  OAI22_X1 U973 ( .A1(n18422), .A2(n18949), .B1(n18958), .B2(n19560), .ZN(
        n3475) );
  OAI22_X1 U974 ( .A1(n18419), .A2(n18949), .B1(n18958), .B2(n19559), .ZN(
        n3459) );
  OAI22_X1 U975 ( .A1(n18440), .A2(n19004), .B1(n19007), .B2(n19558), .ZN(
        n9038) );
  OAI22_X1 U976 ( .A1(n18437), .A2(n19005), .B1(n19007), .B2(n19557), .ZN(
        n9039) );
  OAI22_X1 U977 ( .A1(n18434), .A2(n19004), .B1(n19007), .B2(n19556), .ZN(
        n9040) );
  OAI22_X1 U978 ( .A1(n18431), .A2(n19005), .B1(n19007), .B2(n19555), .ZN(
        n9041) );
  OAI22_X1 U979 ( .A1(n18428), .A2(n19004), .B1(n19006), .B2(n19554), .ZN(
        n9042) );
  OAI22_X1 U980 ( .A1(n18425), .A2(n19005), .B1(n19006), .B2(n19553), .ZN(
        n9043) );
  OAI22_X1 U981 ( .A1(n18422), .A2(n19004), .B1(n19006), .B2(n19552), .ZN(
        n9044) );
  OAI22_X1 U982 ( .A1(n18419), .A2(n19005), .B1(n19006), .B2(n19551), .ZN(
        n9045) );
  OAI22_X1 U983 ( .A1(n18512), .A2(n18950), .B1(n18951), .B2(n19550), .ZN(
        n3955) );
  OAI22_X1 U984 ( .A1(n18509), .A2(n18949), .B1(n18951), .B2(n19549), .ZN(
        n3939) );
  OAI22_X1 U985 ( .A1(n18506), .A2(n18950), .B1(n18951), .B2(n19548), .ZN(
        n3923) );
  OAI22_X1 U986 ( .A1(n18503), .A2(n18949), .B1(n18951), .B2(n19547), .ZN(
        n3907) );
  OAI22_X1 U987 ( .A1(n18500), .A2(n18950), .B1(n18952), .B2(n19546), .ZN(
        n3891) );
  OAI22_X1 U988 ( .A1(n18497), .A2(n18949), .B1(n18952), .B2(n19545), .ZN(
        n3875) );
  OAI22_X1 U989 ( .A1(n18494), .A2(n18950), .B1(n18952), .B2(n19544), .ZN(
        n3859) );
  OAI22_X1 U990 ( .A1(n18491), .A2(n18949), .B1(n18952), .B2(n19543), .ZN(
        n3843) );
  OAI22_X1 U991 ( .A1(n18512), .A2(n18993), .B1(n19002), .B2(n19342), .ZN(
        n8982) );
  OAI22_X1 U992 ( .A1(n18509), .A2(n18993), .B1(n19002), .B2(n19341), .ZN(
        n8983) );
  OAI22_X1 U993 ( .A1(n18506), .A2(n18993), .B1(n19002), .B2(n19340), .ZN(
        n8984) );
  OAI22_X1 U994 ( .A1(n18503), .A2(n18993), .B1(n19002), .B2(n19339), .ZN(
        n8985) );
  OAI22_X1 U995 ( .A1(n18497), .A2(n18993), .B1(n19001), .B2(n19337), .ZN(
        n8987) );
  OAI22_X1 U996 ( .A1(n18494), .A2(n18993), .B1(n19001), .B2(n19336), .ZN(
        n8988) );
  OAI22_X1 U997 ( .A1(n18491), .A2(n18993), .B1(n19001), .B2(n19335), .ZN(
        n8989) );
  OAI22_X1 U998 ( .A1(n18488), .A2(n18993), .B1(n19001), .B2(n19334), .ZN(
        n8990) );
  OAI22_X1 U999 ( .A1(n18485), .A2(n18993), .B1(n19000), .B2(n19333), .ZN(
        n8991) );
  OAI22_X1 U1000 ( .A1(n18482), .A2(n18993), .B1(n19000), .B2(n19332), .ZN(
        n8992) );
  OAI22_X1 U1001 ( .A1(n18479), .A2(n18993), .B1(n19000), .B2(n19331), .ZN(
        n8993) );
  OAI22_X1 U1002 ( .A1(n18476), .A2(n18994), .B1(n19000), .B2(n19330), .ZN(
        n8994) );
  OAI22_X1 U1003 ( .A1(n18473), .A2(n18994), .B1(n18999), .B2(n19329), .ZN(
        n8995) );
  OAI22_X1 U1004 ( .A1(n18470), .A2(n18994), .B1(n18999), .B2(n19328), .ZN(
        n8996) );
  OAI22_X1 U1005 ( .A1(n18467), .A2(n18994), .B1(n18999), .B2(n19327), .ZN(
        n8997) );
  OAI22_X1 U1006 ( .A1(n18461), .A2(n18994), .B1(n18998), .B2(n19325), .ZN(
        n8999) );
  OAI22_X1 U1007 ( .A1(n18455), .A2(n18994), .B1(n18998), .B2(n19323), .ZN(
        n9001) );
  OAI22_X1 U1008 ( .A1(n18449), .A2(n18994), .B1(n18998), .B2(n19321), .ZN(
        n9003) );
  OAI22_X1 U1009 ( .A1(n18446), .A2(n18994), .B1(n18997), .B2(n19320), .ZN(
        n9004) );
  OAI22_X1 U1010 ( .A1(n18443), .A2(n18994), .B1(n18997), .B2(n19319), .ZN(
        n9005) );
  OAI22_X1 U1011 ( .A1(n18488), .A2(n18917), .B1(n18920), .B2(n19318), .ZN(
        n3821) );
  OAI22_X1 U1012 ( .A1(n18485), .A2(n18917), .B1(n18920), .B2(n19317), .ZN(
        n3805) );
  OAI22_X1 U1013 ( .A1(n18482), .A2(n18917), .B1(n18920), .B2(n19316), .ZN(
        n3789) );
  OAI22_X1 U1014 ( .A1(n18479), .A2(n18917), .B1(n18920), .B2(n19315), .ZN(
        n3773) );
  OAI22_X1 U1015 ( .A1(n18476), .A2(n18917), .B1(n18921), .B2(n19314), .ZN(
        n3757) );
  OAI22_X1 U1016 ( .A1(n18473), .A2(n18917), .B1(n18921), .B2(n19313), .ZN(
        n3741) );
  OAI22_X1 U1017 ( .A1(n18470), .A2(n18917), .B1(n18921), .B2(n19312), .ZN(
        n3725) );
  OAI22_X1 U1018 ( .A1(n18467), .A2(n18917), .B1(n18921), .B2(n19311), .ZN(
        n3709) );
  OAI22_X1 U1019 ( .A1(n18464), .A2(n18917), .B1(n18922), .B2(n19310), .ZN(
        n3693) );
  OAI22_X1 U1020 ( .A1(n18461), .A2(n18917), .B1(n18922), .B2(n19309), .ZN(
        n3677) );
  OAI22_X1 U1021 ( .A1(n18458), .A2(n18917), .B1(n18922), .B2(n19308), .ZN(
        n3661) );
  OAI22_X1 U1022 ( .A1(n18455), .A2(n18917), .B1(n18923), .B2(n19307), .ZN(
        n3645) );
  OAI22_X1 U1023 ( .A1(n18449), .A2(n18916), .B1(n18923), .B2(n19305), .ZN(
        n3613) );
  OAI22_X1 U1024 ( .A1(n18446), .A2(n18916), .B1(n18923), .B2(n19304), .ZN(
        n3597) );
  OAI22_X1 U1025 ( .A1(n18443), .A2(n18916), .B1(n18923), .B2(n19303), .ZN(
        n3581) );
  OAI22_X1 U1026 ( .A1(n18440), .A2(n18916), .B1(n18924), .B2(n19302), .ZN(
        n3565) );
  OAI22_X1 U1027 ( .A1(n18437), .A2(n18916), .B1(n18924), .B2(n19301), .ZN(
        n3549) );
  OAI22_X1 U1028 ( .A1(n18434), .A2(n18916), .B1(n18924), .B2(n19300), .ZN(
        n3533) );
  OAI22_X1 U1029 ( .A1(n18431), .A2(n18916), .B1(n18924), .B2(n19299), .ZN(
        n3517) );
  OAI22_X1 U1030 ( .A1(n18428), .A2(n18916), .B1(n18925), .B2(n19298), .ZN(
        n3501) );
  OAI22_X1 U1031 ( .A1(n18425), .A2(n18916), .B1(n18925), .B2(n19297), .ZN(
        n3485) );
  OAI22_X1 U1032 ( .A1(n18422), .A2(n18916), .B1(n18925), .B2(n19296), .ZN(
        n3469) );
  OAI22_X1 U1033 ( .A1(n18419), .A2(n18916), .B1(n18925), .B2(n19295), .ZN(
        n3453) );
  OAI22_X1 U1034 ( .A1(n18440), .A2(n18993), .B1(n18997), .B2(n19214), .ZN(
        n9006) );
  OAI22_X1 U1035 ( .A1(n18437), .A2(n18994), .B1(n18996), .B2(n19213), .ZN(
        n9007) );
  OAI22_X1 U1036 ( .A1(n18434), .A2(n18993), .B1(n18998), .B2(n19212), .ZN(
        n9008) );
  OAI22_X1 U1037 ( .A1(n18431), .A2(n18994), .B1(n18996), .B2(n19211), .ZN(
        n9009) );
  OAI22_X1 U1038 ( .A1(n18428), .A2(n18993), .B1(n18996), .B2(n19210), .ZN(
        n9010) );
  OAI22_X1 U1039 ( .A1(n18425), .A2(n18994), .B1(n18997), .B2(n19209), .ZN(
        n9011) );
  OAI22_X1 U1040 ( .A1(n18422), .A2(n18993), .B1(n18996), .B2(n19208), .ZN(
        n9012) );
  OAI22_X1 U1041 ( .A1(n18419), .A2(n18994), .B1(n18999), .B2(n19207), .ZN(
        n9013) );
  OAI22_X1 U1042 ( .A1(n18512), .A2(n18917), .B1(n18922), .B2(n19206), .ZN(
        n3949) );
  OAI22_X1 U1043 ( .A1(n18509), .A2(n18916), .B1(n18918), .B2(n19205), .ZN(
        n3933) );
  OAI22_X1 U1044 ( .A1(n18506), .A2(n18917), .B1(n18918), .B2(n19204), .ZN(
        n3917) );
  OAI22_X1 U1045 ( .A1(n18503), .A2(n18916), .B1(n18918), .B2(n19203), .ZN(
        n3901) );
  OAI22_X1 U1046 ( .A1(n18500), .A2(n18917), .B1(n18919), .B2(n19202), .ZN(
        n3885) );
  OAI22_X1 U1047 ( .A1(n18497), .A2(n18916), .B1(n18919), .B2(n19201), .ZN(
        n3869) );
  OAI22_X1 U1048 ( .A1(n18494), .A2(n18917), .B1(n18919), .B2(n19200), .ZN(
        n3853) );
  OAI22_X1 U1049 ( .A1(n18491), .A2(n18916), .B1(n18919), .B2(n19199), .ZN(
        n3837) );
  OAI22_X1 U1050 ( .A1(n18490), .A2(n18708), .B1(n18711), .B2(n19166), .ZN(
        n13848) );
  OAI22_X1 U1051 ( .A1(n18487), .A2(n18708), .B1(n18711), .B2(n19165), .ZN(
        n13847) );
  OAI22_X1 U1052 ( .A1(n18484), .A2(n18708), .B1(n18711), .B2(n19164), .ZN(
        n13846) );
  OAI22_X1 U1053 ( .A1(n18481), .A2(n18708), .B1(n18711), .B2(n19163), .ZN(
        n13845) );
  OAI22_X1 U1054 ( .A1(n18478), .A2(n18708), .B1(n18712), .B2(n19162), .ZN(
        n13844) );
  OAI22_X1 U1055 ( .A1(n18475), .A2(n18708), .B1(n18712), .B2(n19161), .ZN(
        n13843) );
  OAI22_X1 U1056 ( .A1(n18472), .A2(n18708), .B1(n18712), .B2(n19160), .ZN(
        n13842) );
  OAI22_X1 U1057 ( .A1(n18469), .A2(n18708), .B1(n18712), .B2(n19159), .ZN(
        n13841) );
  OAI22_X1 U1058 ( .A1(n18466), .A2(n18708), .B1(n18713), .B2(n19158), .ZN(
        n13840) );
  OAI22_X1 U1059 ( .A1(n18463), .A2(n18708), .B1(n18713), .B2(n19157), .ZN(
        n13839) );
  OAI22_X1 U1060 ( .A1(n18460), .A2(n18708), .B1(n18713), .B2(n19156), .ZN(
        n13838) );
  OAI22_X1 U1061 ( .A1(n18457), .A2(n18708), .B1(n18713), .B2(n19155), .ZN(
        n13837) );
  OAI22_X1 U1062 ( .A1(n18454), .A2(n18707), .B1(n18714), .B2(n19154), .ZN(
        n13836) );
  OAI22_X1 U1063 ( .A1(n18451), .A2(n18707), .B1(n18714), .B2(n19153), .ZN(
        n13835) );
  OAI22_X1 U1064 ( .A1(n18448), .A2(n18707), .B1(n18714), .B2(n19152), .ZN(
        n13834) );
  OAI22_X1 U1065 ( .A1(n18445), .A2(n18707), .B1(n18714), .B2(n19151), .ZN(
        n13833) );
  OAI22_X1 U1066 ( .A1(n18442), .A2(n18707), .B1(n18715), .B2(n19150), .ZN(
        n13832) );
  OAI22_X1 U1067 ( .A1(n18439), .A2(n18707), .B1(n18715), .B2(n19149), .ZN(
        n13831) );
  OAI22_X1 U1068 ( .A1(n18436), .A2(n18707), .B1(n18715), .B2(n19148), .ZN(
        n13830) );
  OAI22_X1 U1069 ( .A1(n18433), .A2(n18707), .B1(n18715), .B2(n19147), .ZN(
        n13829) );
  OAI22_X1 U1070 ( .A1(n18430), .A2(n18707), .B1(n18716), .B2(n19146), .ZN(
        n13828) );
  OAI22_X1 U1071 ( .A1(n18427), .A2(n18707), .B1(n18716), .B2(n19145), .ZN(
        n13827) );
  OAI22_X1 U1072 ( .A1(n18424), .A2(n18707), .B1(n18716), .B2(n19144), .ZN(
        n13826) );
  OAI22_X1 U1073 ( .A1(n18421), .A2(n18707), .B1(n18716), .B2(n19143), .ZN(
        n13825) );
  OAI22_X1 U1074 ( .A1(n18514), .A2(n18708), .B1(n18709), .B2(n19134), .ZN(
        n13856) );
  OAI22_X1 U1075 ( .A1(n18511), .A2(n18707), .B1(n18709), .B2(n19133), .ZN(
        n13855) );
  OAI22_X1 U1076 ( .A1(n18508), .A2(n18708), .B1(n18709), .B2(n19132), .ZN(
        n13854) );
  OAI22_X1 U1077 ( .A1(n18505), .A2(n18707), .B1(n18709), .B2(n19131), .ZN(
        n13853) );
  OAI22_X1 U1078 ( .A1(n18502), .A2(n18708), .B1(n18710), .B2(n19130), .ZN(
        n13852) );
  OAI22_X1 U1079 ( .A1(n18499), .A2(n18707), .B1(n18710), .B2(n19129), .ZN(
        n13851) );
  OAI22_X1 U1080 ( .A1(n18496), .A2(n18708), .B1(n18710), .B2(n19128), .ZN(
        n13850) );
  OAI22_X1 U1081 ( .A1(n18493), .A2(n18707), .B1(n18710), .B2(n19127), .ZN(
        n13849) );
  NAND2_X1 U1082 ( .A1(n2199), .A2(n2203), .ZN(n1616) );
  NAND2_X1 U1083 ( .A1(n2198), .A2(n2203), .ZN(n1617) );
  NAND2_X1 U1084 ( .A1(n1584), .A2(n1573), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n1586), .A2(n1579), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n899), .A2(n900), .ZN(n898) );
  NAND2_X1 U1087 ( .A1(n936), .A2(n937), .ZN(n904) );
  NAND2_X1 U1088 ( .A1(n1580), .A2(n1574), .ZN(n987) );
  NAND2_X1 U1089 ( .A1(n1581), .A2(n1574), .ZN(n986) );
  NAND2_X1 U1090 ( .A1(n2210), .A2(n2199), .ZN(n1630) );
  NAND2_X1 U1091 ( .A1(n2210), .A2(n2198), .ZN(n1631) );
  NAND2_X1 U1092 ( .A1(n2213), .A2(n2199), .ZN(n1640) );
  NAND2_X1 U1093 ( .A1(n2213), .A2(n2198), .ZN(n1641) );
  NAND2_X1 U1094 ( .A1(n1586), .A2(n1584), .ZN(n1016) );
  NAND2_X1 U1095 ( .A1(n1583), .A2(n1584), .ZN(n992) );
  NAND2_X1 U1096 ( .A1(n1583), .A2(n1575), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1586), .A2(n1575), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1457), .A2(n1458), .ZN(N696) );
  NOR4_X1 U1099 ( .A1(n1459), .A2(n1460), .A3(n1461), .A4(n1462), .ZN(n1458)
         );
  NOR4_X1 U1100 ( .A1(n1467), .A2(n1468), .A3(n1469), .A4(n1470), .ZN(n1457)
         );
  OAI221_X1 U1101 ( .B1(n19768), .B2(n18668), .C1(n19826), .C2(n18665), .A(
        n1466), .ZN(n1459) );
  NAND2_X1 U1102 ( .A1(n975), .A2(n976), .ZN(N721) );
  NOR4_X1 U1103 ( .A1(n977), .A2(n978), .A3(n979), .A4(n980), .ZN(n976) );
  NOR4_X1 U1104 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n975) );
  OAI221_X1 U1105 ( .B1(n19631), .B2(n18670), .C1(n19655), .C2(n18667), .A(
        n998), .ZN(n977) );
  NAND2_X1 U1106 ( .A1(n1061), .A2(n1062), .ZN(N718) );
  NOR4_X1 U1107 ( .A1(n1063), .A2(n1064), .A3(n1065), .A4(n1066), .ZN(n1062)
         );
  NOR4_X1 U1108 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1061)
         );
  OAI221_X1 U1109 ( .B1(n19634), .B2(n18670), .C1(n19658), .C2(n18667), .A(
        n1070), .ZN(n1063) );
  NAND2_X1 U1110 ( .A1(n1133), .A2(n1134), .ZN(N714) );
  NOR4_X1 U1111 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n1138), .ZN(n1134)
         );
  NOR4_X1 U1112 ( .A1(n1143), .A2(n1144), .A3(n1145), .A4(n1146), .ZN(n1133)
         );
  OAI221_X1 U1113 ( .B1(n19638), .B2(n18670), .C1(n19662), .C2(n18667), .A(
        n1142), .ZN(n1135) );
  NAND2_X1 U1114 ( .A1(n1565), .A2(n1566), .ZN(N690) );
  NOR4_X1 U1115 ( .A1(n1567), .A2(n1568), .A3(n1569), .A4(n1570), .ZN(n1566)
         );
  NOR4_X1 U1116 ( .A1(n1587), .A2(n1588), .A3(n1589), .A4(n1590), .ZN(n1565)
         );
  OAI221_X1 U1117 ( .B1(n19774), .B2(n18668), .C1(n19832), .C2(n18665), .A(
        n1585), .ZN(n1567) );
  NAND2_X1 U1118 ( .A1(n1511), .A2(n1512), .ZN(N693) );
  NOR4_X1 U1119 ( .A1(n1513), .A2(n1514), .A3(n1515), .A4(n1516), .ZN(n1512)
         );
  NOR4_X1 U1120 ( .A1(n1521), .A2(n1522), .A3(n1523), .A4(n1524), .ZN(n1511)
         );
  OAI221_X1 U1121 ( .B1(n19771), .B2(n18668), .C1(n19829), .C2(n18665), .A(
        n1520), .ZN(n1513) );
  NAND2_X1 U1122 ( .A1(n1043), .A2(n1044), .ZN(N719) );
  NOR4_X1 U1123 ( .A1(n1045), .A2(n1046), .A3(n1047), .A4(n1048), .ZN(n1044)
         );
  NOR4_X1 U1124 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1043)
         );
  OAI221_X1 U1125 ( .B1(n19633), .B2(n18670), .C1(n19657), .C2(n18667), .A(
        n1052), .ZN(n1045) );
  NAND2_X1 U1126 ( .A1(n1115), .A2(n1116), .ZN(N715) );
  NOR4_X1 U1127 ( .A1(n1117), .A2(n1118), .A3(n1119), .A4(n1120), .ZN(n1116)
         );
  NOR4_X1 U1128 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1115)
         );
  OAI221_X1 U1129 ( .B1(n19637), .B2(n18670), .C1(n19661), .C2(n18667), .A(
        n1124), .ZN(n1117) );
  NAND2_X1 U1130 ( .A1(n1439), .A2(n1440), .ZN(N697) );
  NOR4_X1 U1131 ( .A1(n1441), .A2(n1442), .A3(n1443), .A4(n1444), .ZN(n1440)
         );
  NOR4_X1 U1132 ( .A1(n1449), .A2(n1450), .A3(n1451), .A4(n1452), .ZN(n1439)
         );
  OAI221_X1 U1133 ( .B1(n19767), .B2(n18668), .C1(n19825), .C2(n18665), .A(
        n1448), .ZN(n1441) );
  NAND2_X1 U1134 ( .A1(n1583), .A2(n1580), .ZN(n1005) );
  NAND2_X1 U1135 ( .A1(n2192), .A2(n2200), .ZN(n1607) );
  NAND2_X1 U1136 ( .A1(n2192), .A2(n2201), .ZN(n1606) );
  NAND2_X1 U1137 ( .A1(n1493), .A2(n1494), .ZN(N694) );
  NOR4_X1 U1138 ( .A1(n1495), .A2(n1496), .A3(n1497), .A4(n1498), .ZN(n1494)
         );
  NOR4_X1 U1139 ( .A1(n1503), .A2(n1504), .A3(n1505), .A4(n1506), .ZN(n1493)
         );
  OAI221_X1 U1140 ( .B1(n19770), .B2(n18668), .C1(n19828), .C2(n18665), .A(
        n1502), .ZN(n1495) );
  NAND2_X1 U1141 ( .A1(n1529), .A2(n1530), .ZN(N692) );
  NOR4_X1 U1142 ( .A1(n1531), .A2(n1532), .A3(n1533), .A4(n1534), .ZN(n1530)
         );
  NOR4_X1 U1143 ( .A1(n1539), .A2(n1540), .A3(n1541), .A4(n1542), .ZN(n1529)
         );
  OAI221_X1 U1144 ( .B1(n19772), .B2(n18668), .C1(n19830), .C2(n18665), .A(
        n1538), .ZN(n1531) );
  NAND2_X1 U1145 ( .A1(n1097), .A2(n1098), .ZN(N716) );
  NOR4_X1 U1146 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1098)
         );
  NOR4_X1 U1147 ( .A1(n1107), .A2(n1108), .A3(n1109), .A4(n1110), .ZN(n1097)
         );
  OAI221_X1 U1148 ( .B1(n19636), .B2(n18670), .C1(n19660), .C2(n18667), .A(
        n1106), .ZN(n1099) );
  NAND2_X1 U1149 ( .A1(n1421), .A2(n1422), .ZN(N698) );
  NOR4_X1 U1150 ( .A1(n1423), .A2(n1424), .A3(n1425), .A4(n1426), .ZN(n1422)
         );
  NOR4_X1 U1151 ( .A1(n1431), .A2(n1432), .A3(n1433), .A4(n1434), .ZN(n1421)
         );
  OAI221_X1 U1152 ( .B1(n19766), .B2(n18668), .C1(n19824), .C2(n18665), .A(
        n1430), .ZN(n1423) );
  NAND2_X1 U1153 ( .A1(n1547), .A2(n1548), .ZN(N691) );
  NOR4_X1 U1154 ( .A1(n1549), .A2(n1550), .A3(n1551), .A4(n1552), .ZN(n1548)
         );
  NOR4_X1 U1155 ( .A1(n1557), .A2(n1558), .A3(n1559), .A4(n1560), .ZN(n1547)
         );
  OAI221_X1 U1156 ( .B1(n19773), .B2(n18668), .C1(n19831), .C2(n18665), .A(
        n1556), .ZN(n1549) );
  NAND2_X1 U1157 ( .A1(n1475), .A2(n1476), .ZN(N695) );
  NOR4_X1 U1158 ( .A1(n1477), .A2(n1478), .A3(n1479), .A4(n1480), .ZN(n1476)
         );
  NOR4_X1 U1159 ( .A1(n1485), .A2(n1486), .A3(n1487), .A4(n1488), .ZN(n1475)
         );
  OAI221_X1 U1160 ( .B1(n19769), .B2(n18668), .C1(n19827), .C2(n18665), .A(
        n1484), .ZN(n1477) );
  NAND2_X1 U1161 ( .A1(n1025), .A2(n1026), .ZN(N720) );
  NOR4_X1 U1162 ( .A1(n1027), .A2(n1028), .A3(n1029), .A4(n1030), .ZN(n1026)
         );
  NOR4_X1 U1163 ( .A1(n1035), .A2(n1036), .A3(n1037), .A4(n1038), .ZN(n1025)
         );
  OAI221_X1 U1164 ( .B1(n19632), .B2(n18670), .C1(n19656), .C2(n18667), .A(
        n1034), .ZN(n1027) );
  NAND2_X1 U1165 ( .A1(n1079), .A2(n1080), .ZN(N717) );
  NOR4_X1 U1166 ( .A1(n1081), .A2(n1082), .A3(n1083), .A4(n1084), .ZN(n1080)
         );
  NOR4_X1 U1167 ( .A1(n1089), .A2(n1090), .A3(n1091), .A4(n1092), .ZN(n1079)
         );
  OAI221_X1 U1168 ( .B1(n19635), .B2(n18670), .C1(n19659), .C2(n18667), .A(
        n1088), .ZN(n1081) );
  NAND2_X1 U1169 ( .A1(n1403), .A2(n1404), .ZN(N699) );
  NOR4_X1 U1170 ( .A1(n1405), .A2(n1406), .A3(n1407), .A4(n1408), .ZN(n1404)
         );
  NOR4_X1 U1171 ( .A1(n1413), .A2(n1414), .A3(n1415), .A4(n1416), .ZN(n1403)
         );
  OAI221_X1 U1172 ( .B1(n19765), .B2(n18668), .C1(n19823), .C2(n18665), .A(
        n1412), .ZN(n1405) );
  AND2_X1 U1173 ( .A1(n1576), .A2(n1573), .ZN(n990) );
  AND2_X1 U1174 ( .A1(n1579), .A2(n1573), .ZN(n989) );
  AND2_X1 U1175 ( .A1(n1577), .A2(n1583), .ZN(n1013) );
  AND2_X1 U1176 ( .A1(n1577), .A2(n1574), .ZN(n1023) );
  NAND2_X1 U1177 ( .A1(n2194), .A2(n2203), .ZN(n1611) );
  NAND2_X1 U1178 ( .A1(n2193), .A2(n2203), .ZN(n1612) );
  AND2_X1 U1179 ( .A1(n1572), .A2(n1583), .ZN(n1014) );
  AND2_X1 U1180 ( .A1(n1572), .A2(n1574), .ZN(n1024) );
  AND2_X1 U1181 ( .A1(n1572), .A2(n1573), .ZN(n985) );
  NAND2_X1 U1182 ( .A1(n2210), .A2(n2194), .ZN(n1625) );
  NAND2_X1 U1183 ( .A1(n2210), .A2(n2193), .ZN(n1626) );
  NAND2_X1 U1184 ( .A1(n2213), .A2(n2194), .ZN(n1635) );
  NAND2_X1 U1185 ( .A1(n2213), .A2(n2193), .ZN(n1636) );
  NAND2_X1 U1186 ( .A1(n2192), .A2(n2196), .ZN(n1601) );
  NAND2_X1 U1187 ( .A1(n2192), .A2(n2195), .ZN(n1602) );
  AND2_X1 U1188 ( .A1(n1583), .A2(n1579), .ZN(n1008) );
  AND2_X1 U1189 ( .A1(n1584), .A2(n1574), .ZN(n1000) );
  AND2_X1 U1190 ( .A1(n1575), .A2(n1573), .ZN(n999) );
  AND2_X1 U1191 ( .A1(n1580), .A2(n1586), .ZN(n1019) );
  AND2_X1 U1192 ( .A1(n1580), .A2(n1573), .ZN(n994) );
  AND2_X1 U1193 ( .A1(n2200), .A2(n2203), .ZN(n1620) );
  AND2_X1 U1194 ( .A1(n2201), .A2(n2203), .ZN(n1619) );
  AND2_X1 U1195 ( .A1(n1581), .A2(n1586), .ZN(n1018) );
  AND2_X1 U1196 ( .A1(n1581), .A2(n1573), .ZN(n995) );
  AND2_X1 U1197 ( .A1(n2192), .A2(n2198), .ZN(n1610) );
  AND2_X1 U1198 ( .A1(n2192), .A2(n2199), .ZN(n1609) );
  AND2_X1 U1199 ( .A1(n1574), .A2(n1575), .ZN(n984) );
  AND2_X1 U1200 ( .A1(n2210), .A2(n2200), .ZN(n1634) );
  AND2_X1 U1201 ( .A1(n2210), .A2(n2201), .ZN(n1633) );
  AND2_X1 U1202 ( .A1(n2213), .A2(n2200), .ZN(n1644) );
  AND2_X1 U1203 ( .A1(n2213), .A2(n2201), .ZN(n1643) );
  AND2_X1 U1204 ( .A1(n1583), .A2(n1581), .ZN(n1009) );
  AND2_X1 U1205 ( .A1(n2192), .A2(n2194), .ZN(n1604) );
  AND2_X1 U1206 ( .A1(n2192), .A2(n2193), .ZN(n1605) );
  AND2_X1 U1207 ( .A1(n2210), .A2(n2196), .ZN(n1628) );
  AND2_X1 U1208 ( .A1(n2210), .A2(n2195), .ZN(n1629) );
  AND2_X1 U1209 ( .A1(n2213), .A2(n2196), .ZN(n1638) );
  AND2_X1 U1210 ( .A1(n2213), .A2(n2195), .ZN(n1639) );
  AND2_X1 U1211 ( .A1(n2196), .A2(n2203), .ZN(n1614) );
  AND2_X1 U1212 ( .A1(n2195), .A2(n2203), .ZN(n1615) );
  INV_X1 U1213 ( .A(DATAIN[8]), .ZN(n19104) );
  INV_X1 U1214 ( .A(DATAIN[31]), .ZN(n19058) );
  INV_X1 U1215 ( .A(DATAIN[3]), .ZN(n19114) );
  INV_X1 U1216 ( .A(DATAIN[4]), .ZN(n19112) );
  INV_X1 U1217 ( .A(DATAIN[5]), .ZN(n19110) );
  INV_X1 U1218 ( .A(DATAIN[6]), .ZN(n19108) );
  INV_X1 U1219 ( .A(DATAIN[7]), .ZN(n19106) );
  INV_X1 U1220 ( .A(DATAIN[9]), .ZN(n19102) );
  INV_X1 U1221 ( .A(DATAIN[10]), .ZN(n19100) );
  INV_X1 U1222 ( .A(DATAIN[11]), .ZN(n19098) );
  INV_X1 U1223 ( .A(DATAIN[12]), .ZN(n19096) );
  INV_X1 U1224 ( .A(DATAIN[13]), .ZN(n19094) );
  INV_X1 U1225 ( .A(DATAIN[14]), .ZN(n19092) );
  INV_X1 U1226 ( .A(DATAIN[15]), .ZN(n19090) );
  INV_X1 U1227 ( .A(DATAIN[16]), .ZN(n19088) );
  INV_X1 U1228 ( .A(DATAIN[17]), .ZN(n19086) );
  INV_X1 U1229 ( .A(DATAIN[18]), .ZN(n19084) );
  INV_X1 U1230 ( .A(DATAIN[19]), .ZN(n19082) );
  INV_X1 U1231 ( .A(DATAIN[20]), .ZN(n19080) );
  INV_X1 U1232 ( .A(DATAIN[21]), .ZN(n19078) );
  INV_X1 U1233 ( .A(DATAIN[22]), .ZN(n19076) );
  INV_X1 U1234 ( .A(DATAIN[23]), .ZN(n19074) );
  INV_X1 U1235 ( .A(DATAIN[24]), .ZN(n19072) );
  INV_X1 U1236 ( .A(DATAIN[25]), .ZN(n19070) );
  INV_X1 U1237 ( .A(DATAIN[26]), .ZN(n19068) );
  INV_X1 U1238 ( .A(DATAIN[27]), .ZN(n19066) );
  INV_X1 U1239 ( .A(DATAIN[28]), .ZN(n19064) );
  INV_X1 U1240 ( .A(DATAIN[29]), .ZN(n19062) );
  INV_X1 U1241 ( .A(DATAIN[30]), .ZN(n19060) );
  INV_X1 U1242 ( .A(DATAIN[0]), .ZN(n19120) );
  INV_X1 U1243 ( .A(DATAIN[1]), .ZN(n19118) );
  INV_X1 U1244 ( .A(DATAIN[2]), .ZN(n19116) );
  NOR3_X1 U1245 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n19124), .ZN(n900) );
  NOR3_X1 U1246 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n19125), .ZN(n937) );
  NOR3_X1 U1247 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n902) );
  NOR3_X1 U1248 ( .A1(n19124), .A2(ADD_WR[1]), .A3(n19126), .ZN(n940) );
  NOR3_X1 U1249 ( .A1(n19124), .A2(ADD_WR[0]), .A3(n19125), .ZN(n959) );
  NOR3_X1 U1250 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n19126), .ZN(n954) );
  NOR3_X1 U1251 ( .A1(n19125), .A2(ADD_WR[2]), .A3(n19126), .ZN(n957) );
  NOR3_X1 U1252 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[2]), .A3(n19921), .ZN(n2199) );
  NOR3_X1 U1253 ( .A1(n19920), .A2(ADD_RD2[2]), .A3(n19921), .ZN(n2198) );
  NOR3_X1 U1254 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[1]), .A3(n19913), .ZN(n1584) );
  NOR3_X1 U1255 ( .A1(n19917), .A2(ADD_RD1[0]), .A3(n19913), .ZN(n1580) );
  NOR3_X1 U1256 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n19920), .ZN(n2200) );
  NOR3_X1 U1257 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(ADD_RD2[0]), .ZN(n2201) );
  NOR3_X1 U1258 ( .A1(n19914), .A2(ADD_RD1[1]), .A3(n19913), .ZN(n1581) );
  AOI22_X1 U1259 ( .A1(n18650), .A2(n17533), .B1(n18649), .B2(n19288), .ZN(
        n1471) );
  NOR4_X1 U1260 ( .A1(n2043), .A2(n2044), .A3(n2045), .A4(n2046), .ZN(n2042)
         );
  OAI221_X1 U1261 ( .B1(n17799), .B2(n18572), .C1(n19766), .C2(n18569), .A(
        n2050), .ZN(n2043) );
  OAI221_X1 U1262 ( .B1(n17903), .B2(n18584), .C1(n17823), .C2(n18581), .A(
        n2049), .ZN(n2044) );
  OAI221_X1 U1263 ( .B1(n19582), .B2(n18596), .C1(n19750), .C2(n18593), .A(
        n2048), .ZN(n2045) );
  NOR4_X1 U1264 ( .A1(n2025), .A2(n2026), .A3(n2027), .A4(n2028), .ZN(n2024)
         );
  OAI221_X1 U1265 ( .B1(n17800), .B2(n18572), .C1(n19765), .C2(n18569), .A(
        n2032), .ZN(n2025) );
  OAI221_X1 U1266 ( .B1(n17904), .B2(n18584), .C1(n17824), .C2(n18581), .A(
        n2031), .ZN(n2026) );
  OAI221_X1 U1267 ( .B1(n19581), .B2(n18596), .C1(n19749), .C2(n18593), .A(
        n2030), .ZN(n2027) );
  NOR4_X1 U1268 ( .A1(n2007), .A2(n2008), .A3(n2009), .A4(n2010), .ZN(n2006)
         );
  OAI221_X1 U1269 ( .B1(n17801), .B2(n18572), .C1(n19764), .C2(n18569), .A(
        n2014), .ZN(n2007) );
  OAI221_X1 U1270 ( .B1(n17905), .B2(n18584), .C1(n17825), .C2(n18581), .A(
        n2013), .ZN(n2008) );
  OAI221_X1 U1271 ( .B1(n19580), .B2(n18596), .C1(n19748), .C2(n18593), .A(
        n2012), .ZN(n2009) );
  NOR4_X1 U1272 ( .A1(n1989), .A2(n1990), .A3(n1991), .A4(n1992), .ZN(n1988)
         );
  OAI221_X1 U1273 ( .B1(n17802), .B2(n18572), .C1(n19763), .C2(n18569), .A(
        n1996), .ZN(n1989) );
  OAI221_X1 U1274 ( .B1(n17906), .B2(n18584), .C1(n17826), .C2(n18581), .A(
        n1995), .ZN(n1990) );
  OAI221_X1 U1275 ( .B1(n19579), .B2(n18596), .C1(n19747), .C2(n18593), .A(
        n1994), .ZN(n1991) );
  NOR4_X1 U1276 ( .A1(n1971), .A2(n1972), .A3(n1973), .A4(n1974), .ZN(n1970)
         );
  OAI221_X1 U1277 ( .B1(n17803), .B2(n18573), .C1(n19762), .C2(n18570), .A(
        n1978), .ZN(n1971) );
  OAI221_X1 U1278 ( .B1(n17907), .B2(n18585), .C1(n17827), .C2(n18582), .A(
        n1977), .ZN(n1972) );
  OAI221_X1 U1279 ( .B1(n19578), .B2(n18597), .C1(n19746), .C2(n18594), .A(
        n1976), .ZN(n1973) );
  NOR4_X1 U1280 ( .A1(n1953), .A2(n1954), .A3(n1955), .A4(n1956), .ZN(n1952)
         );
  OAI221_X1 U1281 ( .B1(n17804), .B2(n18573), .C1(n19761), .C2(n18570), .A(
        n1960), .ZN(n1953) );
  OAI221_X1 U1282 ( .B1(n17908), .B2(n18585), .C1(n17828), .C2(n18582), .A(
        n1959), .ZN(n1954) );
  OAI221_X1 U1283 ( .B1(n19577), .B2(n18597), .C1(n19745), .C2(n18594), .A(
        n1958), .ZN(n1955) );
  NOR4_X1 U1284 ( .A1(n1935), .A2(n1936), .A3(n1937), .A4(n1938), .ZN(n1934)
         );
  OAI221_X1 U1285 ( .B1(n17805), .B2(n18573), .C1(n19760), .C2(n18570), .A(
        n1942), .ZN(n1935) );
  OAI221_X1 U1286 ( .B1(n17909), .B2(n18585), .C1(n17829), .C2(n18582), .A(
        n1941), .ZN(n1936) );
  OAI221_X1 U1287 ( .B1(n19576), .B2(n18597), .C1(n19744), .C2(n18594), .A(
        n1940), .ZN(n1937) );
  NOR4_X1 U1288 ( .A1(n1917), .A2(n1918), .A3(n1919), .A4(n1920), .ZN(n1916)
         );
  OAI221_X1 U1289 ( .B1(n17806), .B2(n18573), .C1(n19759), .C2(n18570), .A(
        n1924), .ZN(n1917) );
  OAI221_X1 U1290 ( .B1(n17910), .B2(n18585), .C1(n17830), .C2(n18582), .A(
        n1923), .ZN(n1918) );
  OAI221_X1 U1291 ( .B1(n19575), .B2(n18597), .C1(n19743), .C2(n18594), .A(
        n1922), .ZN(n1919) );
  NOR4_X1 U1292 ( .A1(n1899), .A2(n1900), .A3(n1901), .A4(n1902), .ZN(n1898)
         );
  OAI221_X1 U1293 ( .B1(n17807), .B2(n18573), .C1(n19758), .C2(n18570), .A(
        n1906), .ZN(n1899) );
  OAI221_X1 U1294 ( .B1(n17911), .B2(n18585), .C1(n17831), .C2(n18582), .A(
        n1905), .ZN(n1900) );
  OAI221_X1 U1295 ( .B1(n19574), .B2(n18597), .C1(n19742), .C2(n18594), .A(
        n1904), .ZN(n1901) );
  NOR4_X1 U1296 ( .A1(n1881), .A2(n1882), .A3(n1883), .A4(n1884), .ZN(n1880)
         );
  OAI221_X1 U1297 ( .B1(n17808), .B2(n18573), .C1(n19757), .C2(n18570), .A(
        n1888), .ZN(n1881) );
  OAI221_X1 U1298 ( .B1(n17912), .B2(n18585), .C1(n17832), .C2(n18582), .A(
        n1887), .ZN(n1882) );
  OAI221_X1 U1299 ( .B1(n19573), .B2(n18597), .C1(n19741), .C2(n18594), .A(
        n1886), .ZN(n1883) );
  NOR4_X1 U1300 ( .A1(n1863), .A2(n1864), .A3(n1865), .A4(n1866), .ZN(n1862)
         );
  OAI221_X1 U1301 ( .B1(n17809), .B2(n18573), .C1(n19756), .C2(n18570), .A(
        n1870), .ZN(n1863) );
  OAI221_X1 U1302 ( .B1(n17913), .B2(n18585), .C1(n17833), .C2(n18582), .A(
        n1869), .ZN(n1864) );
  OAI221_X1 U1303 ( .B1(n19572), .B2(n18597), .C1(n19740), .C2(n18594), .A(
        n1868), .ZN(n1865) );
  NOR4_X1 U1304 ( .A1(n1845), .A2(n1846), .A3(n1847), .A4(n1848), .ZN(n1844)
         );
  OAI221_X1 U1305 ( .B1(n17810), .B2(n18573), .C1(n19755), .C2(n18570), .A(
        n1852), .ZN(n1845) );
  OAI221_X1 U1306 ( .B1(n17914), .B2(n18585), .C1(n17834), .C2(n18582), .A(
        n1851), .ZN(n1846) );
  OAI221_X1 U1307 ( .B1(n19571), .B2(n18597), .C1(n19739), .C2(n18594), .A(
        n1850), .ZN(n1847) );
  NOR4_X1 U1308 ( .A1(n1827), .A2(n1828), .A3(n1829), .A4(n1830), .ZN(n1826)
         );
  OAI221_X1 U1309 ( .B1(n17811), .B2(n18573), .C1(n19754), .C2(n18570), .A(
        n1834), .ZN(n1827) );
  OAI221_X1 U1310 ( .B1(n17915), .B2(n18585), .C1(n17835), .C2(n18582), .A(
        n1833), .ZN(n1828) );
  OAI221_X1 U1311 ( .B1(n19570), .B2(n18597), .C1(n19738), .C2(n18594), .A(
        n1832), .ZN(n1829) );
  NOR4_X1 U1312 ( .A1(n1809), .A2(n1810), .A3(n1811), .A4(n1812), .ZN(n1808)
         );
  OAI221_X1 U1313 ( .B1(n17812), .B2(n18573), .C1(n19753), .C2(n18570), .A(
        n1816), .ZN(n1809) );
  OAI221_X1 U1314 ( .B1(n17916), .B2(n18585), .C1(n17836), .C2(n18582), .A(
        n1815), .ZN(n1810) );
  OAI221_X1 U1315 ( .B1(n19569), .B2(n18597), .C1(n19737), .C2(n18594), .A(
        n1814), .ZN(n1811) );
  NOR4_X1 U1316 ( .A1(n1791), .A2(n1792), .A3(n1793), .A4(n1794), .ZN(n1790)
         );
  OAI221_X1 U1317 ( .B1(n17813), .B2(n18573), .C1(n19752), .C2(n18570), .A(
        n1798), .ZN(n1791) );
  OAI221_X1 U1318 ( .B1(n17917), .B2(n18585), .C1(n17837), .C2(n18582), .A(
        n1797), .ZN(n1792) );
  OAI221_X1 U1319 ( .B1(n19568), .B2(n18597), .C1(n19736), .C2(n18594), .A(
        n1796), .ZN(n1793) );
  NOR4_X1 U1320 ( .A1(n1773), .A2(n1774), .A3(n1775), .A4(n1776), .ZN(n1772)
         );
  OAI221_X1 U1321 ( .B1(n17814), .B2(n18573), .C1(n19751), .C2(n18570), .A(
        n1780), .ZN(n1773) );
  OAI221_X1 U1322 ( .B1(n17918), .B2(n18585), .C1(n17838), .C2(n18582), .A(
        n1779), .ZN(n1774) );
  OAI221_X1 U1323 ( .B1(n19567), .B2(n18597), .C1(n19735), .C2(n18594), .A(
        n1778), .ZN(n1775) );
  NOR4_X1 U1324 ( .A1(n1755), .A2(n1756), .A3(n1757), .A4(n1758), .ZN(n1754)
         );
  OAI221_X1 U1325 ( .B1(n18195), .B2(n18574), .C1(n19638), .C2(n18571), .A(
        n1762), .ZN(n1755) );
  OAI221_X1 U1326 ( .B1(n18227), .B2(n18586), .C1(n18203), .C2(n18583), .A(
        n1761), .ZN(n1756) );
  OAI221_X1 U1327 ( .B1(n19566), .B2(n18598), .C1(n19734), .C2(n18595), .A(
        n1760), .ZN(n1757) );
  NOR4_X1 U1328 ( .A1(n1737), .A2(n1738), .A3(n1739), .A4(n1740), .ZN(n1736)
         );
  OAI221_X1 U1329 ( .B1(n18196), .B2(n18574), .C1(n19637), .C2(n18571), .A(
        n1744), .ZN(n1737) );
  OAI221_X1 U1330 ( .B1(n18228), .B2(n18586), .C1(n18204), .C2(n18583), .A(
        n1743), .ZN(n1738) );
  OAI221_X1 U1331 ( .B1(n19565), .B2(n18598), .C1(n19733), .C2(n18595), .A(
        n1742), .ZN(n1739) );
  NOR4_X1 U1332 ( .A1(n1719), .A2(n1720), .A3(n1721), .A4(n1722), .ZN(n1718)
         );
  OAI221_X1 U1333 ( .B1(n18197), .B2(n18574), .C1(n19636), .C2(n18571), .A(
        n1726), .ZN(n1719) );
  OAI221_X1 U1334 ( .B1(n18229), .B2(n18586), .C1(n18205), .C2(n18583), .A(
        n1725), .ZN(n1720) );
  OAI221_X1 U1335 ( .B1(n19564), .B2(n18598), .C1(n19732), .C2(n18595), .A(
        n1724), .ZN(n1721) );
  NOR4_X1 U1336 ( .A1(n1701), .A2(n1702), .A3(n1703), .A4(n1704), .ZN(n1700)
         );
  OAI221_X1 U1337 ( .B1(n18198), .B2(n18574), .C1(n19635), .C2(n18571), .A(
        n1708), .ZN(n1701) );
  OAI221_X1 U1338 ( .B1(n18230), .B2(n18586), .C1(n18206), .C2(n18583), .A(
        n1707), .ZN(n1702) );
  OAI221_X1 U1339 ( .B1(n19563), .B2(n18598), .C1(n19731), .C2(n18595), .A(
        n1706), .ZN(n1703) );
  NOR4_X1 U1340 ( .A1(n1683), .A2(n1684), .A3(n1685), .A4(n1686), .ZN(n1682)
         );
  OAI221_X1 U1341 ( .B1(n18199), .B2(n18574), .C1(n19634), .C2(n18571), .A(
        n1690), .ZN(n1683) );
  OAI221_X1 U1342 ( .B1(n18231), .B2(n18586), .C1(n18207), .C2(n18583), .A(
        n1689), .ZN(n1684) );
  OAI221_X1 U1343 ( .B1(n19562), .B2(n18598), .C1(n19730), .C2(n18595), .A(
        n1688), .ZN(n1685) );
  NOR4_X1 U1344 ( .A1(n1665), .A2(n1666), .A3(n1667), .A4(n1668), .ZN(n1664)
         );
  OAI221_X1 U1345 ( .B1(n18200), .B2(n18574), .C1(n19633), .C2(n18571), .A(
        n1672), .ZN(n1665) );
  OAI221_X1 U1346 ( .B1(n18232), .B2(n18586), .C1(n18208), .C2(n18583), .A(
        n1671), .ZN(n1666) );
  OAI221_X1 U1347 ( .B1(n19561), .B2(n18598), .C1(n19729), .C2(n18595), .A(
        n1670), .ZN(n1667) );
  NOR4_X1 U1348 ( .A1(n1647), .A2(n1648), .A3(n1649), .A4(n1650), .ZN(n1646)
         );
  OAI221_X1 U1349 ( .B1(n18201), .B2(n18574), .C1(n19632), .C2(n18571), .A(
        n1654), .ZN(n1647) );
  OAI221_X1 U1350 ( .B1(n18233), .B2(n18586), .C1(n18209), .C2(n18583), .A(
        n1653), .ZN(n1648) );
  OAI221_X1 U1351 ( .B1(n19560), .B2(n18598), .C1(n19728), .C2(n18595), .A(
        n1652), .ZN(n1649) );
  NOR4_X1 U1352 ( .A1(n1597), .A2(n1598), .A3(n1599), .A4(n1600), .ZN(n1596)
         );
  OAI221_X1 U1353 ( .B1(n18202), .B2(n18574), .C1(n19631), .C2(n18571), .A(
        n1618), .ZN(n1597) );
  OAI221_X1 U1354 ( .B1(n18234), .B2(n18586), .C1(n18210), .C2(n18583), .A(
        n1613), .ZN(n1598) );
  OAI221_X1 U1355 ( .B1(n19559), .B2(n18598), .C1(n19727), .C2(n18595), .A(
        n1608), .ZN(n1599) );
  NOR4_X1 U1356 ( .A1(n2205), .A2(n2206), .A3(n2207), .A4(n2208), .ZN(n2185)
         );
  OAI221_X1 U1357 ( .B1(n18099), .B2(n18524), .C1(n19832), .C2(n18521), .A(
        n2214), .ZN(n2205) );
  OAI221_X1 U1358 ( .B1(n19726), .B2(n18548), .C1(n19822), .C2(n18545), .A(
        n2211), .ZN(n2207) );
  OAI221_X1 U1359 ( .B1(n17847), .B2(n18536), .C1(n18123), .C2(n18533), .A(
        n2212), .ZN(n2206) );
  NOR4_X1 U1360 ( .A1(n2177), .A2(n2178), .A3(n2179), .A4(n2180), .ZN(n2167)
         );
  OAI221_X1 U1361 ( .B1(n18100), .B2(n18524), .C1(n19831), .C2(n18521), .A(
        n2184), .ZN(n2177) );
  OAI221_X1 U1362 ( .B1(n19725), .B2(n18548), .C1(n19821), .C2(n18545), .A(
        n2182), .ZN(n2179) );
  OAI221_X1 U1363 ( .B1(n17848), .B2(n18536), .C1(n18124), .C2(n18533), .A(
        n2183), .ZN(n2178) );
  NOR4_X1 U1364 ( .A1(n2159), .A2(n2160), .A3(n2161), .A4(n2162), .ZN(n2149)
         );
  OAI221_X1 U1365 ( .B1(n18101), .B2(n18524), .C1(n19830), .C2(n18521), .A(
        n2166), .ZN(n2159) );
  OAI221_X1 U1366 ( .B1(n19724), .B2(n18548), .C1(n19820), .C2(n18545), .A(
        n2164), .ZN(n2161) );
  OAI221_X1 U1367 ( .B1(n17849), .B2(n18536), .C1(n18125), .C2(n18533), .A(
        n2165), .ZN(n2160) );
  NOR4_X1 U1368 ( .A1(n2141), .A2(n2142), .A3(n2143), .A4(n2144), .ZN(n2131)
         );
  OAI221_X1 U1369 ( .B1(n18102), .B2(n18524), .C1(n19829), .C2(n18521), .A(
        n2148), .ZN(n2141) );
  OAI221_X1 U1370 ( .B1(n19723), .B2(n18548), .C1(n19819), .C2(n18545), .A(
        n2146), .ZN(n2143) );
  OAI221_X1 U1371 ( .B1(n17850), .B2(n18536), .C1(n18126), .C2(n18533), .A(
        n2147), .ZN(n2142) );
  NOR4_X1 U1372 ( .A1(n2123), .A2(n2124), .A3(n2125), .A4(n2126), .ZN(n2113)
         );
  OAI221_X1 U1373 ( .B1(n18103), .B2(n18524), .C1(n19828), .C2(n18521), .A(
        n2130), .ZN(n2123) );
  OAI221_X1 U1374 ( .B1(n19722), .B2(n18548), .C1(n19818), .C2(n18545), .A(
        n2128), .ZN(n2125) );
  OAI221_X1 U1375 ( .B1(n17851), .B2(n18536), .C1(n18127), .C2(n18533), .A(
        n2129), .ZN(n2124) );
  NOR4_X1 U1376 ( .A1(n2105), .A2(n2106), .A3(n2107), .A4(n2108), .ZN(n2095)
         );
  OAI221_X1 U1377 ( .B1(n18104), .B2(n18524), .C1(n19827), .C2(n18521), .A(
        n2112), .ZN(n2105) );
  OAI221_X1 U1378 ( .B1(n19721), .B2(n18548), .C1(n19817), .C2(n18545), .A(
        n2110), .ZN(n2107) );
  OAI221_X1 U1379 ( .B1(n17852), .B2(n18536), .C1(n18128), .C2(n18533), .A(
        n2111), .ZN(n2106) );
  NOR4_X1 U1380 ( .A1(n2087), .A2(n2088), .A3(n2089), .A4(n2090), .ZN(n2077)
         );
  OAI221_X1 U1381 ( .B1(n18105), .B2(n18524), .C1(n19826), .C2(n18521), .A(
        n2094), .ZN(n2087) );
  OAI221_X1 U1382 ( .B1(n19720), .B2(n18548), .C1(n19816), .C2(n18545), .A(
        n2092), .ZN(n2089) );
  OAI221_X1 U1383 ( .B1(n17853), .B2(n18536), .C1(n18129), .C2(n18533), .A(
        n2093), .ZN(n2088) );
  NOR4_X1 U1384 ( .A1(n2069), .A2(n2070), .A3(n2071), .A4(n2072), .ZN(n2059)
         );
  OAI221_X1 U1385 ( .B1(n18106), .B2(n18524), .C1(n19825), .C2(n18521), .A(
        n2076), .ZN(n2069) );
  OAI221_X1 U1386 ( .B1(n19719), .B2(n18548), .C1(n19815), .C2(n18545), .A(
        n2074), .ZN(n2071) );
  OAI221_X1 U1387 ( .B1(n17854), .B2(n18536), .C1(n18130), .C2(n18533), .A(
        n2075), .ZN(n2070) );
  AND3_X1 U1388 ( .A1(n970), .A2(n19123), .A3(ADD_WR[4]), .ZN(n899) );
  AND3_X1 U1389 ( .A1(ADD_WR[4]), .A2(n970), .A3(ADD_WR[3]), .ZN(n936) );
  AND3_X1 U1390 ( .A1(n970), .A2(n19122), .A3(ADD_WR[3]), .ZN(n939) );
  OAI221_X1 U1391 ( .B1(n17871), .B2(n18656), .C1(n18171), .C2(n18653), .A(
        n1591), .ZN(n1590) );
  AOI22_X1 U1392 ( .A1(n18650), .A2(n17527), .B1(n18649), .B2(n19294), .ZN(
        n1591) );
  OAI221_X1 U1393 ( .B1(n17881), .B2(n18656), .C1(n18181), .C2(n18653), .A(
        n1399), .ZN(n1398) );
  AOI22_X1 U1394 ( .A1(n18650), .A2(n17537), .B1(n18648), .B2(n19284), .ZN(
        n1399) );
  OAI221_X1 U1395 ( .B1(n17882), .B2(n18656), .C1(n18182), .C2(n18653), .A(
        n1381), .ZN(n1380) );
  AOI22_X1 U1396 ( .A1(n18650), .A2(n17538), .B1(n18648), .B2(n19283), .ZN(
        n1381) );
  OAI221_X1 U1397 ( .B1(n17883), .B2(n18657), .C1(n18183), .C2(n18654), .A(
        n1363), .ZN(n1362) );
  AOI22_X1 U1398 ( .A1(n18651), .A2(n17539), .B1(n18648), .B2(n19282), .ZN(
        n1363) );
  OAI221_X1 U1399 ( .B1(n17888), .B2(n18657), .C1(n18188), .C2(n18654), .A(
        n1273), .ZN(n1272) );
  AOI22_X1 U1400 ( .A1(n18651), .A2(n17544), .B1(n18648), .B2(n19277), .ZN(
        n1273) );
  OAI221_X1 U1401 ( .B1(n17889), .B2(n18657), .C1(n18189), .C2(n18654), .A(
        n1255), .ZN(n1254) );
  AOI22_X1 U1402 ( .A1(n18651), .A2(n17545), .B1(n18648), .B2(n19276), .ZN(
        n1255) );
  OAI221_X1 U1403 ( .B1(n17890), .B2(n18657), .C1(n18190), .C2(n18654), .A(
        n1237), .ZN(n1236) );
  AOI22_X1 U1404 ( .A1(n18651), .A2(n17546), .B1(n18648), .B2(n19275), .ZN(
        n1237) );
  OAI221_X1 U1405 ( .B1(n17872), .B2(n18656), .C1(n18172), .C2(n18653), .A(
        n1561), .ZN(n1560) );
  AOI22_X1 U1406 ( .A1(n18650), .A2(n17528), .B1(n18649), .B2(n19293), .ZN(
        n1561) );
  OAI221_X1 U1407 ( .B1(n17884), .B2(n18657), .C1(n18184), .C2(n18654), .A(
        n1345), .ZN(n1344) );
  AOI22_X1 U1408 ( .A1(n18651), .A2(n17540), .B1(n18648), .B2(n19281), .ZN(
        n1345) );
  OAI221_X1 U1409 ( .B1(n17885), .B2(n18657), .C1(n18185), .C2(n18654), .A(
        n1327), .ZN(n1326) );
  AOI22_X1 U1410 ( .A1(n18651), .A2(n17541), .B1(n18648), .B2(n19280), .ZN(
        n1327) );
  OAI221_X1 U1411 ( .B1(n17886), .B2(n18657), .C1(n18186), .C2(n18654), .A(
        n1309), .ZN(n1308) );
  AOI22_X1 U1412 ( .A1(n18651), .A2(n17542), .B1(n18648), .B2(n19279), .ZN(
        n1309) );
  OAI221_X1 U1413 ( .B1(n17887), .B2(n18657), .C1(n18187), .C2(n18654), .A(
        n1291), .ZN(n1290) );
  AOI22_X1 U1414 ( .A1(n18651), .A2(n17543), .B1(n18648), .B2(n19278), .ZN(
        n1291) );
  OAI221_X1 U1415 ( .B1(n17891), .B2(n18657), .C1(n18191), .C2(n18654), .A(
        n1219), .ZN(n1218) );
  AOI22_X1 U1416 ( .A1(n18651), .A2(n17547), .B1(n18647), .B2(n19274), .ZN(
        n1219) );
  OAI221_X1 U1417 ( .B1(n17892), .B2(n18657), .C1(n18192), .C2(n18654), .A(
        n1201), .ZN(n1200) );
  AOI22_X1 U1418 ( .A1(n18651), .A2(n17548), .B1(n18647), .B2(n19273), .ZN(
        n1201) );
  OAI221_X1 U1419 ( .B1(n17893), .B2(n18657), .C1(n18193), .C2(n18654), .A(
        n1183), .ZN(n1182) );
  AOI22_X1 U1420 ( .A1(n18651), .A2(n17549), .B1(n18647), .B2(n19272), .ZN(
        n1183) );
  OAI221_X1 U1421 ( .B1(n17894), .B2(n18657), .C1(n18194), .C2(n18654), .A(
        n1165), .ZN(n1164) );
  AOI22_X1 U1422 ( .A1(n18651), .A2(n17550), .B1(n18647), .B2(n19271), .ZN(
        n1165) );
  OAI221_X1 U1423 ( .B1(n17878), .B2(n18656), .C1(n18178), .C2(n18653), .A(
        n1453), .ZN(n1452) );
  AOI22_X1 U1424 ( .A1(n18650), .A2(n17534), .B1(n18649), .B2(n19287), .ZN(
        n1453) );
  OAI221_X1 U1425 ( .B1(n17879), .B2(n18656), .C1(n18179), .C2(n18653), .A(
        n1435), .ZN(n1434) );
  AOI22_X1 U1426 ( .A1(n18650), .A2(n17535), .B1(n18648), .B2(n19286), .ZN(
        n1435) );
  OAI221_X1 U1427 ( .B1(n17880), .B2(n18656), .C1(n18180), .C2(n18653), .A(
        n1417), .ZN(n1416) );
  AOI22_X1 U1428 ( .A1(n18650), .A2(n17536), .B1(n18648), .B2(n19285), .ZN(
        n1417) );
  OAI221_X1 U1429 ( .B1(n17874), .B2(n18656), .C1(n18174), .C2(n18653), .A(
        n1525), .ZN(n1524) );
  AOI22_X1 U1430 ( .A1(n18650), .A2(n17530), .B1(n18649), .B2(n19291), .ZN(
        n1525) );
  OAI221_X1 U1431 ( .B1(n18226), .B2(n18658), .C1(n18322), .C2(n18655), .A(
        n1007), .ZN(n1004) );
  AOI22_X1 U1432 ( .A1(n18652), .A2(n17670), .B1(n18647), .B2(n19191), .ZN(
        n1007) );
  OAI221_X1 U1433 ( .B1(n17875), .B2(n18656), .C1(n18175), .C2(n18653), .A(
        n1507), .ZN(n1506) );
  AOI22_X1 U1434 ( .A1(n18650), .A2(n17531), .B1(n18649), .B2(n19290), .ZN(
        n1507) );
  OAI221_X1 U1435 ( .B1(n17876), .B2(n18656), .C1(n18176), .C2(n18653), .A(
        n1489), .ZN(n1488) );
  AOI22_X1 U1436 ( .A1(n18650), .A2(n17532), .B1(n18649), .B2(n19289), .ZN(
        n1489) );
  OAI221_X1 U1437 ( .B1(n18223), .B2(n18658), .C1(n18319), .C2(n18655), .A(
        n1075), .ZN(n1074) );
  AOI22_X1 U1438 ( .A1(n18652), .A2(n17667), .B1(n18647), .B2(n19194), .ZN(
        n1075) );
  OAI221_X1 U1439 ( .B1(n18224), .B2(n18658), .C1(n18320), .C2(n18655), .A(
        n1057), .ZN(n1056) );
  AOI22_X1 U1440 ( .A1(n18652), .A2(n17668), .B1(n18647), .B2(n19193), .ZN(
        n1057) );
  OAI221_X1 U1441 ( .B1(n17873), .B2(n18656), .C1(n18173), .C2(n18653), .A(
        n1543), .ZN(n1542) );
  AOI22_X1 U1442 ( .A1(n18650), .A2(n17529), .B1(n18649), .B2(n19292), .ZN(
        n1543) );
  OAI221_X1 U1443 ( .B1(n18225), .B2(n18658), .C1(n18321), .C2(n18655), .A(
        n1039), .ZN(n1038) );
  AOI22_X1 U1444 ( .A1(n18652), .A2(n17669), .B1(n18647), .B2(n19192), .ZN(
        n1039) );
  OAI221_X1 U1445 ( .B1(n18219), .B2(n18658), .C1(n18315), .C2(n18655), .A(
        n1147), .ZN(n1146) );
  AOI22_X1 U1446 ( .A1(n18652), .A2(n17663), .B1(n18647), .B2(n19198), .ZN(
        n1147) );
  OAI221_X1 U1447 ( .B1(n18220), .B2(n18658), .C1(n18316), .C2(n18655), .A(
        n1129), .ZN(n1128) );
  AOI22_X1 U1448 ( .A1(n18652), .A2(n17664), .B1(n18647), .B2(n19197), .ZN(
        n1129) );
  OAI221_X1 U1449 ( .B1(n18221), .B2(n18658), .C1(n18317), .C2(n18655), .A(
        n1111), .ZN(n1110) );
  AOI22_X1 U1450 ( .A1(n18652), .A2(n17665), .B1(n18647), .B2(n19196), .ZN(
        n1111) );
  OAI221_X1 U1451 ( .B1(n18222), .B2(n18658), .C1(n18318), .C2(n18655), .A(
        n1093), .ZN(n1092) );
  AOI22_X1 U1452 ( .A1(n18652), .A2(n17666), .B1(n18647), .B2(n19195), .ZN(
        n1093) );
  OAI221_X1 U1453 ( .B1(n17871), .B2(n18560), .C1(n18171), .C2(n18557), .A(
        n2209), .ZN(n2208) );
  AOI22_X1 U1454 ( .A1(n18554), .A2(n18275), .B1(n18553), .B2(n19294), .ZN(
        n2209) );
  OAI221_X1 U1455 ( .B1(n17872), .B2(n18560), .C1(n18172), .C2(n18557), .A(
        n2181), .ZN(n2180) );
  AOI22_X1 U1456 ( .A1(n18554), .A2(n18276), .B1(n18553), .B2(n19293), .ZN(
        n2181) );
  OAI221_X1 U1457 ( .B1(n17873), .B2(n18560), .C1(n18173), .C2(n18557), .A(
        n2163), .ZN(n2162) );
  AOI22_X1 U1458 ( .A1(n18554), .A2(n18277), .B1(n18553), .B2(n19292), .ZN(
        n2163) );
  OAI221_X1 U1459 ( .B1(n17874), .B2(n18560), .C1(n18174), .C2(n18557), .A(
        n2145), .ZN(n2144) );
  AOI22_X1 U1460 ( .A1(n18554), .A2(n18278), .B1(n18553), .B2(n19291), .ZN(
        n2145) );
  OAI221_X1 U1461 ( .B1(n17875), .B2(n18560), .C1(n18175), .C2(n18557), .A(
        n2127), .ZN(n2126) );
  AOI22_X1 U1462 ( .A1(n18554), .A2(n18279), .B1(n18553), .B2(n19290), .ZN(
        n2127) );
  OAI221_X1 U1463 ( .B1(n17876), .B2(n18560), .C1(n18176), .C2(n18557), .A(
        n2109), .ZN(n2108) );
  AOI22_X1 U1464 ( .A1(n18554), .A2(n18280), .B1(n18553), .B2(n19289), .ZN(
        n2109) );
  OAI221_X1 U1465 ( .B1(n17878), .B2(n18560), .C1(n18178), .C2(n18557), .A(
        n2073), .ZN(n2072) );
  AOI22_X1 U1466 ( .A1(n18554), .A2(n18282), .B1(n18553), .B2(n19287), .ZN(
        n2073) );
  OAI221_X1 U1467 ( .B1(n18091), .B2(n18610), .C1(n19840), .C2(n18607), .A(
        n1759), .ZN(n1758) );
  AOI22_X1 U1468 ( .A1(n18604), .A2(n19246), .B1(n18599), .B2(n19896), .ZN(
        n1759) );
  OAI221_X1 U1469 ( .B1(n18219), .B2(n18562), .C1(n18315), .C2(n18559), .A(
        n1767), .ZN(n1766) );
  AOI22_X1 U1470 ( .A1(n18556), .A2(n18067), .B1(n18551), .B2(n19198), .ZN(
        n1767) );
  OAI221_X1 U1471 ( .B1(n18092), .B2(n18610), .C1(n19839), .C2(n18607), .A(
        n1741), .ZN(n1740) );
  AOI22_X1 U1472 ( .A1(n18604), .A2(n19245), .B1(n18599), .B2(n19895), .ZN(
        n1741) );
  OAI221_X1 U1473 ( .B1(n18220), .B2(n18562), .C1(n18316), .C2(n18559), .A(
        n1749), .ZN(n1748) );
  AOI22_X1 U1474 ( .A1(n18556), .A2(n18068), .B1(n18551), .B2(n19197), .ZN(
        n1749) );
  OAI221_X1 U1475 ( .B1(n18093), .B2(n18610), .C1(n19838), .C2(n18607), .A(
        n1723), .ZN(n1722) );
  AOI22_X1 U1476 ( .A1(n18604), .A2(n19244), .B1(n18599), .B2(n19894), .ZN(
        n1723) );
  OAI221_X1 U1477 ( .B1(n18221), .B2(n18562), .C1(n18317), .C2(n18559), .A(
        n1731), .ZN(n1730) );
  AOI22_X1 U1478 ( .A1(n18556), .A2(n18069), .B1(n18551), .B2(n19196), .ZN(
        n1731) );
  OAI221_X1 U1479 ( .B1(n18094), .B2(n18610), .C1(n19837), .C2(n18607), .A(
        n1705), .ZN(n1704) );
  AOI22_X1 U1480 ( .A1(n18604), .A2(n19243), .B1(n18599), .B2(n19893), .ZN(
        n1705) );
  OAI221_X1 U1481 ( .B1(n18222), .B2(n18562), .C1(n18318), .C2(n18559), .A(
        n1713), .ZN(n1712) );
  AOI22_X1 U1482 ( .A1(n18556), .A2(n18070), .B1(n18551), .B2(n19195), .ZN(
        n1713) );
  OAI221_X1 U1483 ( .B1(n18095), .B2(n18610), .C1(n19836), .C2(n18607), .A(
        n1687), .ZN(n1686) );
  AOI22_X1 U1484 ( .A1(n18604), .A2(n19242), .B1(n18599), .B2(n19892), .ZN(
        n1687) );
  OAI221_X1 U1485 ( .B1(n18223), .B2(n18562), .C1(n18319), .C2(n18559), .A(
        n1695), .ZN(n1694) );
  AOI22_X1 U1486 ( .A1(n18556), .A2(n18071), .B1(n18551), .B2(n19194), .ZN(
        n1695) );
  OAI221_X1 U1487 ( .B1(n18096), .B2(n18610), .C1(n19835), .C2(n18607), .A(
        n1669), .ZN(n1668) );
  AOI22_X1 U1488 ( .A1(n18604), .A2(n19241), .B1(n18599), .B2(n19891), .ZN(
        n1669) );
  OAI221_X1 U1489 ( .B1(n18224), .B2(n18562), .C1(n18320), .C2(n18559), .A(
        n1677), .ZN(n1676) );
  AOI22_X1 U1490 ( .A1(n18556), .A2(n18072), .B1(n18551), .B2(n19193), .ZN(
        n1677) );
  OAI221_X1 U1491 ( .B1(n18097), .B2(n18610), .C1(n19834), .C2(n18607), .A(
        n1651), .ZN(n1650) );
  AOI22_X1 U1492 ( .A1(n18604), .A2(n19240), .B1(n18599), .B2(n19890), .ZN(
        n1651) );
  OAI221_X1 U1493 ( .B1(n18225), .B2(n18562), .C1(n18321), .C2(n18559), .A(
        n1659), .ZN(n1658) );
  AOI22_X1 U1494 ( .A1(n18556), .A2(n18073), .B1(n18551), .B2(n19192), .ZN(
        n1659) );
  OAI221_X1 U1495 ( .B1(n18098), .B2(n18610), .C1(n19833), .C2(n18607), .A(
        n1603), .ZN(n1600) );
  AOI22_X1 U1496 ( .A1(n18604), .A2(n19239), .B1(n18599), .B2(n19889), .ZN(
        n1603) );
  OAI221_X1 U1497 ( .B1(n18226), .B2(n18562), .C1(n18322), .C2(n18559), .A(
        n1627), .ZN(n1624) );
  AOI22_X1 U1498 ( .A1(n18556), .A2(n18074), .B1(n18551), .B2(n19191), .ZN(
        n1627) );
  OAI221_X1 U1499 ( .B1(n19727), .B2(n18706), .C1(n2215), .C2(n18703), .A(n983), .ZN(n980) );
  AOI22_X1 U1500 ( .A1(n18700), .A2(n19255), .B1(n18695), .B2(n17622), .ZN(
        n983) );
  OAI221_X1 U1501 ( .B1(n19730), .B2(n18706), .C1(n2242), .C2(n18703), .A(
        n1067), .ZN(n1066) );
  AOI22_X1 U1502 ( .A1(n18700), .A2(n19258), .B1(n18695), .B2(n17619), .ZN(
        n1067) );
  OAI221_X1 U1503 ( .B1(n19729), .B2(n18706), .C1(n2233), .C2(n18703), .A(
        n1049), .ZN(n1048) );
  AOI22_X1 U1504 ( .A1(n18700), .A2(n19257), .B1(n18695), .B2(n17620), .ZN(
        n1049) );
  OAI221_X1 U1505 ( .B1(n19728), .B2(n18706), .C1(n2224), .C2(n18703), .A(
        n1031), .ZN(n1030) );
  AOI22_X1 U1506 ( .A1(n18700), .A2(n19256), .B1(n18695), .B2(n17621), .ZN(
        n1031) );
  OAI221_X1 U1507 ( .B1(n19734), .B2(n18706), .C1(n2278), .C2(n18703), .A(
        n1139), .ZN(n1138) );
  AOI22_X1 U1508 ( .A1(n18700), .A2(n19262), .B1(n18695), .B2(n17615), .ZN(
        n1139) );
  OAI221_X1 U1509 ( .B1(n19733), .B2(n18706), .C1(n2269), .C2(n18703), .A(
        n1121), .ZN(n1120) );
  AOI22_X1 U1510 ( .A1(n18700), .A2(n19261), .B1(n18695), .B2(n17616), .ZN(
        n1121) );
  OAI221_X1 U1511 ( .B1(n19732), .B2(n18706), .C1(n2260), .C2(n18703), .A(
        n1103), .ZN(n1102) );
  AOI22_X1 U1512 ( .A1(n18700), .A2(n19260), .B1(n18695), .B2(n17617), .ZN(
        n1103) );
  OAI221_X1 U1513 ( .B1(n19731), .B2(n18706), .C1(n2251), .C2(n18703), .A(
        n1085), .ZN(n1084) );
  AOI22_X1 U1514 ( .A1(n18700), .A2(n19259), .B1(n18695), .B2(n17618), .ZN(
        n1085) );
  OAI221_X1 U1515 ( .B1(n17877), .B2(n18560), .C1(n18177), .C2(n18557), .A(
        n2091), .ZN(n2090) );
  AOI22_X1 U1516 ( .A1(n18554), .A2(n18281), .B1(n18553), .B2(n19288), .ZN(
        n2091) );
  OAI221_X1 U1517 ( .B1(n19630), .B2(n18704), .C1(n2494), .C2(n18701), .A(
        n1571), .ZN(n1570) );
  AOI22_X1 U1518 ( .A1(n18698), .A2(n19494), .B1(n18697), .B2(n17687), .ZN(
        n1571) );
  OAI221_X1 U1519 ( .B1(n19748), .B2(n18704), .C1(n2404), .C2(n18701), .A(
        n1391), .ZN(n1390) );
  AOI22_X1 U1520 ( .A1(n18698), .A2(n19484), .B1(n18696), .B2(n17601), .ZN(
        n1391) );
  OAI221_X1 U1521 ( .B1(n19747), .B2(n18704), .C1(n2395), .C2(n18701), .A(
        n1373), .ZN(n1372) );
  AOI22_X1 U1522 ( .A1(n18698), .A2(n19483), .B1(n18696), .B2(n17602), .ZN(
        n1373) );
  OAI221_X1 U1523 ( .B1(n19746), .B2(n18705), .C1(n2386), .C2(n18702), .A(
        n1355), .ZN(n1354) );
  AOI22_X1 U1524 ( .A1(n18699), .A2(n19482), .B1(n18696), .B2(n17603), .ZN(
        n1355) );
  OAI221_X1 U1525 ( .B1(n19741), .B2(n18705), .C1(n2341), .C2(n18702), .A(
        n1265), .ZN(n1264) );
  AOI22_X1 U1526 ( .A1(n18699), .A2(n19477), .B1(n18696), .B2(n17608), .ZN(
        n1265) );
  OAI221_X1 U1527 ( .B1(n19740), .B2(n18705), .C1(n2332), .C2(n18702), .A(
        n1247), .ZN(n1246) );
  AOI22_X1 U1528 ( .A1(n18699), .A2(n19476), .B1(n18696), .B2(n17609), .ZN(
        n1247) );
  OAI221_X1 U1529 ( .B1(n19739), .B2(n18705), .C1(n2323), .C2(n18702), .A(
        n1229), .ZN(n1228) );
  AOI22_X1 U1530 ( .A1(n18699), .A2(n19475), .B1(n18696), .B2(n17610), .ZN(
        n1229) );
  OAI221_X1 U1531 ( .B1(n19629), .B2(n18704), .C1(n2485), .C2(n18701), .A(
        n1553), .ZN(n1552) );
  AOI22_X1 U1532 ( .A1(n18698), .A2(n19493), .B1(n18697), .B2(n17688), .ZN(
        n1553) );
  OAI221_X1 U1533 ( .B1(n19745), .B2(n18705), .C1(n2377), .C2(n18702), .A(
        n1337), .ZN(n1336) );
  AOI22_X1 U1534 ( .A1(n18699), .A2(n19481), .B1(n18696), .B2(n17604), .ZN(
        n1337) );
  OAI221_X1 U1535 ( .B1(n19744), .B2(n18705), .C1(n2368), .C2(n18702), .A(
        n1319), .ZN(n1318) );
  AOI22_X1 U1536 ( .A1(n18699), .A2(n19480), .B1(n18696), .B2(n17605), .ZN(
        n1319) );
  OAI221_X1 U1537 ( .B1(n19743), .B2(n18705), .C1(n2359), .C2(n18702), .A(
        n1301), .ZN(n1300) );
  AOI22_X1 U1538 ( .A1(n18699), .A2(n19479), .B1(n18696), .B2(n17606), .ZN(
        n1301) );
  OAI221_X1 U1539 ( .B1(n19742), .B2(n18705), .C1(n2350), .C2(n18702), .A(
        n1283), .ZN(n1282) );
  AOI22_X1 U1540 ( .A1(n18699), .A2(n19478), .B1(n18696), .B2(n17607), .ZN(
        n1283) );
  OAI221_X1 U1541 ( .B1(n19738), .B2(n18705), .C1(n2314), .C2(n18702), .A(
        n1211), .ZN(n1210) );
  AOI22_X1 U1542 ( .A1(n18699), .A2(n19474), .B1(n18695), .B2(n17611), .ZN(
        n1211) );
  OAI221_X1 U1543 ( .B1(n19737), .B2(n18705), .C1(n2305), .C2(n18702), .A(
        n1193), .ZN(n1192) );
  AOI22_X1 U1544 ( .A1(n18699), .A2(n19473), .B1(n18695), .B2(n17612), .ZN(
        n1193) );
  OAI221_X1 U1545 ( .B1(n19736), .B2(n18705), .C1(n2296), .C2(n18702), .A(
        n1175), .ZN(n1174) );
  AOI22_X1 U1546 ( .A1(n18699), .A2(n19472), .B1(n18695), .B2(n17613), .ZN(
        n1175) );
  OAI221_X1 U1547 ( .B1(n19735), .B2(n18705), .C1(n2287), .C2(n18702), .A(
        n1157), .ZN(n1156) );
  AOI22_X1 U1548 ( .A1(n18699), .A2(n19471), .B1(n18695), .B2(n17614), .ZN(
        n1157) );
  OAI221_X1 U1549 ( .B1(n19624), .B2(n18704), .C1(n2440), .C2(n18701), .A(
        n1463), .ZN(n1462) );
  AOI22_X1 U1550 ( .A1(n18698), .A2(n19488), .B1(n18697), .B2(n17693), .ZN(
        n1463) );
  OAI221_X1 U1551 ( .B1(n19623), .B2(n18704), .C1(n2431), .C2(n18701), .A(
        n1445), .ZN(n1444) );
  AOI22_X1 U1552 ( .A1(n18698), .A2(n19487), .B1(n18697), .B2(n17694), .ZN(
        n1445) );
  OAI221_X1 U1553 ( .B1(n19750), .B2(n18704), .C1(n2422), .C2(n18701), .A(
        n1427), .ZN(n1426) );
  AOI22_X1 U1554 ( .A1(n18698), .A2(n19486), .B1(n18696), .B2(n17599), .ZN(
        n1427) );
  OAI221_X1 U1555 ( .B1(n19749), .B2(n18704), .C1(n2413), .C2(n18701), .A(
        n1409), .ZN(n1408) );
  AOI22_X1 U1556 ( .A1(n18698), .A2(n19485), .B1(n18696), .B2(n17600), .ZN(
        n1409) );
  OAI221_X1 U1557 ( .B1(n19627), .B2(n18704), .C1(n2467), .C2(n18701), .A(
        n1517), .ZN(n1516) );
  AOI22_X1 U1558 ( .A1(n18698), .A2(n19491), .B1(n18697), .B2(n17690), .ZN(
        n1517) );
  OAI221_X1 U1559 ( .B1(n19626), .B2(n18704), .C1(n2458), .C2(n18701), .A(
        n1499), .ZN(n1498) );
  AOI22_X1 U1560 ( .A1(n18698), .A2(n19490), .B1(n18697), .B2(n17691), .ZN(
        n1499) );
  OAI221_X1 U1561 ( .B1(n19625), .B2(n18704), .C1(n2449), .C2(n18701), .A(
        n1481), .ZN(n1480) );
  AOI22_X1 U1562 ( .A1(n18698), .A2(n19489), .B1(n18697), .B2(n17692), .ZN(
        n1481) );
  OAI221_X1 U1563 ( .B1(n19628), .B2(n18704), .C1(n2476), .C2(n18701), .A(
        n1535), .ZN(n1534) );
  AOI22_X1 U1564 ( .A1(n18698), .A2(n19492), .B1(n18697), .B2(n17689), .ZN(
        n1535) );
  OAI221_X1 U1565 ( .B1(n18123), .B2(n18644), .C1(n19606), .C2(n18641), .A(
        n1592), .ZN(n1589) );
  AOI22_X1 U1566 ( .A1(n18638), .A2(n19230), .B1(n18637), .B2(n17575), .ZN(
        n1592) );
  OAI221_X1 U1567 ( .B1(n18133), .B2(n18644), .C1(n19596), .C2(n18641), .A(
        n1400), .ZN(n1397) );
  AOI22_X1 U1568 ( .A1(n18638), .A2(n19388), .B1(n18636), .B2(n17585), .ZN(
        n1400) );
  OAI221_X1 U1569 ( .B1(n18134), .B2(n18644), .C1(n19595), .C2(n18641), .A(
        n1382), .ZN(n1379) );
  AOI22_X1 U1570 ( .A1(n18638), .A2(n19387), .B1(n18636), .B2(n17586), .ZN(
        n1382) );
  OAI221_X1 U1571 ( .B1(n18135), .B2(n18645), .C1(n19594), .C2(n18642), .A(
        n1364), .ZN(n1361) );
  AOI22_X1 U1572 ( .A1(n18639), .A2(n19386), .B1(n18636), .B2(n17587), .ZN(
        n1364) );
  OAI221_X1 U1573 ( .B1(n18140), .B2(n18645), .C1(n19589), .C2(n18642), .A(
        n1274), .ZN(n1271) );
  AOI22_X1 U1574 ( .A1(n18639), .A2(n19381), .B1(n18636), .B2(n17592), .ZN(
        n1274) );
  OAI221_X1 U1575 ( .B1(n18141), .B2(n18645), .C1(n19588), .C2(n18642), .A(
        n1256), .ZN(n1253) );
  AOI22_X1 U1576 ( .A1(n18639), .A2(n19380), .B1(n18636), .B2(n17593), .ZN(
        n1256) );
  OAI221_X1 U1577 ( .B1(n18142), .B2(n18645), .C1(n19587), .C2(n18642), .A(
        n1238), .ZN(n1235) );
  AOI22_X1 U1578 ( .A1(n18639), .A2(n19379), .B1(n18636), .B2(n17594), .ZN(
        n1238) );
  OAI221_X1 U1579 ( .B1(n18124), .B2(n18644), .C1(n19605), .C2(n18641), .A(
        n1562), .ZN(n1559) );
  AOI22_X1 U1580 ( .A1(n18638), .A2(n19229), .B1(n18637), .B2(n17576), .ZN(
        n1562) );
  OAI221_X1 U1581 ( .B1(n18136), .B2(n18645), .C1(n19593), .C2(n18642), .A(
        n1346), .ZN(n1343) );
  AOI22_X1 U1582 ( .A1(n18639), .A2(n19385), .B1(n18636), .B2(n17588), .ZN(
        n1346) );
  OAI221_X1 U1583 ( .B1(n18137), .B2(n18645), .C1(n19592), .C2(n18642), .A(
        n1328), .ZN(n1325) );
  AOI22_X1 U1584 ( .A1(n18639), .A2(n19384), .B1(n18636), .B2(n17589), .ZN(
        n1328) );
  OAI221_X1 U1585 ( .B1(n18138), .B2(n18645), .C1(n19591), .C2(n18642), .A(
        n1310), .ZN(n1307) );
  AOI22_X1 U1586 ( .A1(n18639), .A2(n19383), .B1(n18636), .B2(n17590), .ZN(
        n1310) );
  OAI221_X1 U1587 ( .B1(n18139), .B2(n18645), .C1(n19590), .C2(n18642), .A(
        n1292), .ZN(n1289) );
  AOI22_X1 U1588 ( .A1(n18639), .A2(n19382), .B1(n18636), .B2(n17591), .ZN(
        n1292) );
  OAI221_X1 U1589 ( .B1(n18143), .B2(n18645), .C1(n19586), .C2(n18642), .A(
        n1220), .ZN(n1217) );
  AOI22_X1 U1590 ( .A1(n18639), .A2(n19378), .B1(n18635), .B2(n17595), .ZN(
        n1220) );
  OAI221_X1 U1591 ( .B1(n18144), .B2(n18645), .C1(n19585), .C2(n18642), .A(
        n1202), .ZN(n1199) );
  AOI22_X1 U1592 ( .A1(n18639), .A2(n19377), .B1(n18635), .B2(n17596), .ZN(
        n1202) );
  OAI221_X1 U1593 ( .B1(n18145), .B2(n18645), .C1(n19584), .C2(n18642), .A(
        n1184), .ZN(n1181) );
  AOI22_X1 U1594 ( .A1(n18639), .A2(n19376), .B1(n18635), .B2(n17597), .ZN(
        n1184) );
  OAI221_X1 U1595 ( .B1(n18146), .B2(n18645), .C1(n19583), .C2(n18642), .A(
        n1166), .ZN(n1163) );
  AOI22_X1 U1596 ( .A1(n18639), .A2(n19375), .B1(n18635), .B2(n17598), .ZN(
        n1166) );
  OAI221_X1 U1597 ( .B1(n18129), .B2(n18644), .C1(n19600), .C2(n18641), .A(
        n1472), .ZN(n1469) );
  AOI22_X1 U1598 ( .A1(n18638), .A2(n19224), .B1(n18637), .B2(n17581), .ZN(
        n1472) );
  OAI221_X1 U1599 ( .B1(n18130), .B2(n18644), .C1(n19599), .C2(n18641), .A(
        n1454), .ZN(n1451) );
  AOI22_X1 U1600 ( .A1(n18638), .A2(n19223), .B1(n18637), .B2(n17582), .ZN(
        n1454) );
  OAI221_X1 U1601 ( .B1(n18131), .B2(n18644), .C1(n19598), .C2(n18641), .A(
        n1436), .ZN(n1433) );
  AOI22_X1 U1602 ( .A1(n18638), .A2(n19390), .B1(n18636), .B2(n17583), .ZN(
        n1436) );
  OAI221_X1 U1603 ( .B1(n18132), .B2(n18644), .C1(n19597), .C2(n18641), .A(
        n1418), .ZN(n1415) );
  AOI22_X1 U1604 ( .A1(n18638), .A2(n19389), .B1(n18636), .B2(n17584), .ZN(
        n1418) );
  OAI221_X1 U1605 ( .B1(n18126), .B2(n18644), .C1(n19603), .C2(n18641), .A(
        n1526), .ZN(n1523) );
  AOI22_X1 U1606 ( .A1(n18638), .A2(n19227), .B1(n18637), .B2(n17578), .ZN(
        n1526) );
  OAI221_X1 U1607 ( .B1(n18306), .B2(n18646), .C1(n19551), .C2(n18643), .A(
        n1012), .ZN(n1003) );
  AOI22_X1 U1608 ( .A1(n18640), .A2(n19367), .B1(n18635), .B2(n17686), .ZN(
        n1012) );
  OAI221_X1 U1609 ( .B1(n18127), .B2(n18644), .C1(n19602), .C2(n18641), .A(
        n1508), .ZN(n1505) );
  AOI22_X1 U1610 ( .A1(n18638), .A2(n19226), .B1(n18637), .B2(n17579), .ZN(
        n1508) );
  OAI221_X1 U1611 ( .B1(n18128), .B2(n18644), .C1(n19601), .C2(n18641), .A(
        n1490), .ZN(n1487) );
  AOI22_X1 U1612 ( .A1(n18638), .A2(n19225), .B1(n18637), .B2(n17580), .ZN(
        n1490) );
  OAI221_X1 U1613 ( .B1(n18303), .B2(n18646), .C1(n19554), .C2(n18643), .A(
        n1076), .ZN(n1073) );
  AOI22_X1 U1614 ( .A1(n18640), .A2(n19370), .B1(n18635), .B2(n17683), .ZN(
        n1076) );
  OAI221_X1 U1615 ( .B1(n18304), .B2(n18646), .C1(n19553), .C2(n18643), .A(
        n1058), .ZN(n1055) );
  AOI22_X1 U1616 ( .A1(n18640), .A2(n19369), .B1(n18635), .B2(n17684), .ZN(
        n1058) );
  OAI221_X1 U1617 ( .B1(n18125), .B2(n18644), .C1(n19604), .C2(n18641), .A(
        n1544), .ZN(n1541) );
  AOI22_X1 U1618 ( .A1(n18638), .A2(n19228), .B1(n18637), .B2(n17577), .ZN(
        n1544) );
  OAI221_X1 U1619 ( .B1(n18305), .B2(n18646), .C1(n19552), .C2(n18643), .A(
        n1040), .ZN(n1037) );
  AOI22_X1 U1620 ( .A1(n18640), .A2(n19368), .B1(n18635), .B2(n17685), .ZN(
        n1040) );
  OAI221_X1 U1621 ( .B1(n18299), .B2(n18646), .C1(n19558), .C2(n18643), .A(
        n1148), .ZN(n1145) );
  AOI22_X1 U1622 ( .A1(n18640), .A2(n19374), .B1(n18635), .B2(n17679), .ZN(
        n1148) );
  OAI221_X1 U1623 ( .B1(n18300), .B2(n18646), .C1(n19557), .C2(n18643), .A(
        n1130), .ZN(n1127) );
  AOI22_X1 U1624 ( .A1(n18640), .A2(n19373), .B1(n18635), .B2(n17680), .ZN(
        n1130) );
  OAI221_X1 U1625 ( .B1(n18301), .B2(n18646), .C1(n19556), .C2(n18643), .A(
        n1112), .ZN(n1109) );
  AOI22_X1 U1626 ( .A1(n18640), .A2(n19372), .B1(n18635), .B2(n17681), .ZN(
        n1112) );
  OAI221_X1 U1627 ( .B1(n18302), .B2(n18646), .C1(n19555), .C2(n18643), .A(
        n1094), .ZN(n1091) );
  AOI22_X1 U1628 ( .A1(n18640), .A2(n19371), .B1(n18635), .B2(n17682), .ZN(
        n1094) );
  OAI221_X1 U1629 ( .B1(n19857), .B2(n18694), .C1(n18234), .C2(n18691), .A(
        n988), .ZN(n979) );
  AOI22_X1 U1630 ( .A1(n18688), .A2(n19215), .B1(n18683), .B2(n17750), .ZN(
        n988) );
  OAI221_X1 U1631 ( .B1(n19860), .B2(n18694), .C1(n18231), .C2(n18691), .A(
        n1068), .ZN(n1065) );
  AOI22_X1 U1632 ( .A1(n18688), .A2(n19218), .B1(n18683), .B2(n17747), .ZN(
        n1068) );
  OAI221_X1 U1633 ( .B1(n19859), .B2(n18694), .C1(n18232), .C2(n18691), .A(
        n1050), .ZN(n1047) );
  AOI22_X1 U1634 ( .A1(n18688), .A2(n19217), .B1(n18683), .B2(n17748), .ZN(
        n1050) );
  OAI221_X1 U1635 ( .B1(n19858), .B2(n18694), .C1(n18233), .C2(n18691), .A(
        n1032), .ZN(n1029) );
  AOI22_X1 U1636 ( .A1(n18688), .A2(n19216), .B1(n18683), .B2(n17749), .ZN(
        n1032) );
  OAI221_X1 U1637 ( .B1(n19864), .B2(n18694), .C1(n18227), .C2(n18691), .A(
        n1140), .ZN(n1137) );
  AOI22_X1 U1638 ( .A1(n18688), .A2(n19222), .B1(n18683), .B2(n17743), .ZN(
        n1140) );
  OAI221_X1 U1639 ( .B1(n19863), .B2(n18694), .C1(n18228), .C2(n18691), .A(
        n1122), .ZN(n1119) );
  AOI22_X1 U1640 ( .A1(n18688), .A2(n19221), .B1(n18683), .B2(n17744), .ZN(
        n1122) );
  OAI221_X1 U1641 ( .B1(n19862), .B2(n18694), .C1(n18229), .C2(n18691), .A(
        n1104), .ZN(n1101) );
  AOI22_X1 U1642 ( .A1(n18688), .A2(n19220), .B1(n18683), .B2(n17745), .ZN(
        n1104) );
  OAI221_X1 U1643 ( .B1(n19861), .B2(n18694), .C1(n18230), .C2(n18691), .A(
        n1086), .ZN(n1083) );
  AOI22_X1 U1644 ( .A1(n18688), .A2(n19219), .B1(n18683), .B2(n17746), .ZN(
        n1086) );
  OAI221_X1 U1645 ( .B1(n19678), .B2(n18692), .C1(n17895), .C2(n18689), .A(
        n1578), .ZN(n1569) );
  AOI22_X1 U1646 ( .A1(n18686), .A2(n19366), .B1(n18685), .B2(n17759), .ZN(
        n1578) );
  OAI221_X1 U1647 ( .B1(n19878), .B2(n18692), .C1(n17905), .C2(n18689), .A(
        n1392), .ZN(n1389) );
  AOI22_X1 U1648 ( .A1(n18686), .A2(n19356), .B1(n18684), .B2(n17729), .ZN(
        n1392) );
  OAI221_X1 U1649 ( .B1(n19877), .B2(n18692), .C1(n17906), .C2(n18689), .A(
        n1374), .ZN(n1371) );
  AOI22_X1 U1650 ( .A1(n18686), .A2(n19355), .B1(n18684), .B2(n17730), .ZN(
        n1374) );
  OAI221_X1 U1651 ( .B1(n19876), .B2(n18693), .C1(n17907), .C2(n18690), .A(
        n1356), .ZN(n1353) );
  AOI22_X1 U1652 ( .A1(n18687), .A2(n19354), .B1(n18684), .B2(n17731), .ZN(
        n1356) );
  OAI221_X1 U1653 ( .B1(n19871), .B2(n18693), .C1(n17912), .C2(n18690), .A(
        n1266), .ZN(n1263) );
  AOI22_X1 U1654 ( .A1(n18687), .A2(n19349), .B1(n18684), .B2(n17736), .ZN(
        n1266) );
  OAI221_X1 U1655 ( .B1(n19870), .B2(n18693), .C1(n17913), .C2(n18690), .A(
        n1248), .ZN(n1245) );
  AOI22_X1 U1656 ( .A1(n18687), .A2(n19348), .B1(n18684), .B2(n17737), .ZN(
        n1248) );
  OAI221_X1 U1657 ( .B1(n19869), .B2(n18693), .C1(n17914), .C2(n18690), .A(
        n1230), .ZN(n1227) );
  AOI22_X1 U1658 ( .A1(n18687), .A2(n19347), .B1(n18684), .B2(n17738), .ZN(
        n1230) );
  OAI221_X1 U1659 ( .B1(n19677), .B2(n18692), .C1(n17896), .C2(n18689), .A(
        n1554), .ZN(n1551) );
  AOI22_X1 U1660 ( .A1(n18686), .A2(n19365), .B1(n18685), .B2(n17760), .ZN(
        n1554) );
  OAI221_X1 U1661 ( .B1(n19875), .B2(n18693), .C1(n17908), .C2(n18690), .A(
        n1338), .ZN(n1335) );
  AOI22_X1 U1662 ( .A1(n18687), .A2(n19353), .B1(n18684), .B2(n17732), .ZN(
        n1338) );
  OAI221_X1 U1663 ( .B1(n19874), .B2(n18693), .C1(n17909), .C2(n18690), .A(
        n1320), .ZN(n1317) );
  AOI22_X1 U1664 ( .A1(n18687), .A2(n19352), .B1(n18684), .B2(n17733), .ZN(
        n1320) );
  OAI221_X1 U1665 ( .B1(n19873), .B2(n18693), .C1(n17910), .C2(n18690), .A(
        n1302), .ZN(n1299) );
  AOI22_X1 U1666 ( .A1(n18687), .A2(n19351), .B1(n18684), .B2(n17734), .ZN(
        n1302) );
  OAI221_X1 U1667 ( .B1(n19872), .B2(n18693), .C1(n17911), .C2(n18690), .A(
        n1284), .ZN(n1281) );
  AOI22_X1 U1668 ( .A1(n18687), .A2(n19350), .B1(n18684), .B2(n17735), .ZN(
        n1284) );
  OAI221_X1 U1669 ( .B1(n19868), .B2(n18693), .C1(n17915), .C2(n18690), .A(
        n1212), .ZN(n1209) );
  AOI22_X1 U1670 ( .A1(n18687), .A2(n19346), .B1(n18683), .B2(n17739), .ZN(
        n1212) );
  OAI221_X1 U1671 ( .B1(n19867), .B2(n18693), .C1(n17916), .C2(n18690), .A(
        n1194), .ZN(n1191) );
  AOI22_X1 U1672 ( .A1(n18687), .A2(n19345), .B1(n18683), .B2(n17740), .ZN(
        n1194) );
  OAI221_X1 U1673 ( .B1(n19866), .B2(n18693), .C1(n17917), .C2(n18690), .A(
        n1176), .ZN(n1173) );
  AOI22_X1 U1674 ( .A1(n18687), .A2(n19344), .B1(n18683), .B2(n17741), .ZN(
        n1176) );
  OAI221_X1 U1675 ( .B1(n19865), .B2(n18693), .C1(n17918), .C2(n18690), .A(
        n1158), .ZN(n1155) );
  AOI22_X1 U1676 ( .A1(n18687), .A2(n19343), .B1(n18683), .B2(n17742), .ZN(
        n1158) );
  OAI221_X1 U1677 ( .B1(n19672), .B2(n18692), .C1(n17901), .C2(n18689), .A(
        n1464), .ZN(n1461) );
  AOI22_X1 U1678 ( .A1(n18686), .A2(n19360), .B1(n18685), .B2(n17765), .ZN(
        n1464) );
  OAI221_X1 U1679 ( .B1(n19671), .B2(n18692), .C1(n17902), .C2(n18689), .A(
        n1446), .ZN(n1443) );
  AOI22_X1 U1680 ( .A1(n18686), .A2(n19359), .B1(n18685), .B2(n17766), .ZN(
        n1446) );
  OAI221_X1 U1681 ( .B1(n19880), .B2(n18692), .C1(n17903), .C2(n18689), .A(
        n1428), .ZN(n1425) );
  AOI22_X1 U1682 ( .A1(n18686), .A2(n19358), .B1(n18684), .B2(n17727), .ZN(
        n1428) );
  OAI221_X1 U1683 ( .B1(n19879), .B2(n18692), .C1(n17904), .C2(n18689), .A(
        n1410), .ZN(n1407) );
  AOI22_X1 U1684 ( .A1(n18686), .A2(n19357), .B1(n18684), .B2(n17728), .ZN(
        n1410) );
  OAI221_X1 U1685 ( .B1(n19675), .B2(n18692), .C1(n17898), .C2(n18689), .A(
        n1518), .ZN(n1515) );
  AOI22_X1 U1686 ( .A1(n18686), .A2(n19363), .B1(n18685), .B2(n17762), .ZN(
        n1518) );
  OAI221_X1 U1687 ( .B1(n19674), .B2(n18692), .C1(n17899), .C2(n18689), .A(
        n1500), .ZN(n1497) );
  AOI22_X1 U1688 ( .A1(n18686), .A2(n19362), .B1(n18685), .B2(n17763), .ZN(
        n1500) );
  OAI221_X1 U1689 ( .B1(n19673), .B2(n18692), .C1(n17900), .C2(n18689), .A(
        n1482), .ZN(n1479) );
  AOI22_X1 U1690 ( .A1(n18686), .A2(n19361), .B1(n18685), .B2(n17764), .ZN(
        n1482) );
  OAI221_X1 U1691 ( .B1(n19676), .B2(n18692), .C1(n17897), .C2(n18689), .A(
        n1536), .ZN(n1533) );
  AOI22_X1 U1692 ( .A1(n18686), .A2(n19364), .B1(n18685), .B2(n17761), .ZN(
        n1536) );
  OAI221_X1 U1693 ( .B1(n18099), .B2(n18632), .C1(n19342), .C2(n18629), .A(
        n1593), .ZN(n1588) );
  AOI22_X1 U1694 ( .A1(n18626), .A2(n19614), .B1(n18625), .B2(n19462), .ZN(
        n1593) );
  OAI221_X1 U1695 ( .B1(n18283), .B2(n18680), .C1(n19206), .C2(n18677), .A(
        n1582), .ZN(n1568) );
  AOI22_X1 U1696 ( .A1(n18674), .A2(n19438), .B1(n18673), .B2(n17655), .ZN(
        n1582) );
  OAI221_X1 U1697 ( .B1(n18109), .B2(n18632), .C1(n19332), .C2(n18629), .A(
        n1401), .ZN(n1396) );
  AOI22_X1 U1698 ( .A1(n18626), .A2(n19700), .B1(n18624), .B2(n19452), .ZN(
        n1401) );
  OAI221_X1 U1699 ( .B1(n18077), .B2(n18680), .C1(n19316), .C2(n18677), .A(
        n1393), .ZN(n1388) );
  AOI22_X1 U1700 ( .A1(n18674), .A2(n19428), .B1(n18672), .B2(n17505), .ZN(
        n1393) );
  OAI221_X1 U1701 ( .B1(n18110), .B2(n18632), .C1(n19331), .C2(n18629), .A(
        n1383), .ZN(n1378) );
  AOI22_X1 U1702 ( .A1(n18626), .A2(n19699), .B1(n18624), .B2(n19451), .ZN(
        n1383) );
  OAI221_X1 U1703 ( .B1(n18078), .B2(n18680), .C1(n19315), .C2(n18677), .A(
        n1375), .ZN(n1370) );
  AOI22_X1 U1704 ( .A1(n18674), .A2(n19427), .B1(n18672), .B2(n17506), .ZN(
        n1375) );
  OAI221_X1 U1705 ( .B1(n18111), .B2(n18633), .C1(n19330), .C2(n18630), .A(
        n1365), .ZN(n1360) );
  AOI22_X1 U1706 ( .A1(n18627), .A2(n19698), .B1(n18624), .B2(n19450), .ZN(
        n1365) );
  OAI221_X1 U1707 ( .B1(n18079), .B2(n18681), .C1(n19314), .C2(n18678), .A(
        n1357), .ZN(n1352) );
  AOI22_X1 U1708 ( .A1(n18675), .A2(n19426), .B1(n18672), .B2(n17507), .ZN(
        n1357) );
  OAI221_X1 U1709 ( .B1(n18116), .B2(n18633), .C1(n19325), .C2(n18630), .A(
        n1275), .ZN(n1270) );
  AOI22_X1 U1710 ( .A1(n18627), .A2(n19693), .B1(n18624), .B2(n19445), .ZN(
        n1275) );
  OAI221_X1 U1711 ( .B1(n18084), .B2(n18681), .C1(n19309), .C2(n18678), .A(
        n1267), .ZN(n1262) );
  AOI22_X1 U1712 ( .A1(n18675), .A2(n19421), .B1(n18672), .B2(n17512), .ZN(
        n1267) );
  OAI221_X1 U1713 ( .B1(n18117), .B2(n18633), .C1(n18045), .C2(n18630), .A(
        n1257), .ZN(n1252) );
  AOI22_X1 U1714 ( .A1(n18627), .A2(n19692), .B1(n18624), .B2(n19444), .ZN(
        n1257) );
  OAI221_X1 U1715 ( .B1(n18085), .B2(n18681), .C1(n19308), .C2(n18678), .A(
        n1249), .ZN(n1244) );
  AOI22_X1 U1716 ( .A1(n18675), .A2(n19420), .B1(n18672), .B2(n17513), .ZN(
        n1249) );
  OAI221_X1 U1717 ( .B1(n18118), .B2(n18633), .C1(n19323), .C2(n18630), .A(
        n1239), .ZN(n1234) );
  AOI22_X1 U1718 ( .A1(n18627), .A2(n19691), .B1(n18624), .B2(n19443), .ZN(
        n1239) );
  OAI221_X1 U1719 ( .B1(n18086), .B2(n18681), .C1(n19307), .C2(n18678), .A(
        n1231), .ZN(n1226) );
  AOI22_X1 U1720 ( .A1(n18675), .A2(n19419), .B1(n18672), .B2(n17514), .ZN(
        n1231) );
  OAI221_X1 U1721 ( .B1(n18100), .B2(n18632), .C1(n19341), .C2(n18629), .A(
        n1563), .ZN(n1558) );
  AOI22_X1 U1722 ( .A1(n18626), .A2(n19613), .B1(n18625), .B2(n19461), .ZN(
        n1563) );
  OAI221_X1 U1723 ( .B1(n18284), .B2(n18680), .C1(n19205), .C2(n18677), .A(
        n1555), .ZN(n1550) );
  AOI22_X1 U1724 ( .A1(n18674), .A2(n19437), .B1(n18673), .B2(n17656), .ZN(
        n1555) );
  OAI221_X1 U1725 ( .B1(n18112), .B2(n18633), .C1(n19329), .C2(n18630), .A(
        n1347), .ZN(n1342) );
  AOI22_X1 U1726 ( .A1(n18627), .A2(n19697), .B1(n18624), .B2(n19449), .ZN(
        n1347) );
  OAI221_X1 U1727 ( .B1(n18080), .B2(n18681), .C1(n19313), .C2(n18678), .A(
        n1339), .ZN(n1334) );
  AOI22_X1 U1728 ( .A1(n18675), .A2(n19425), .B1(n18672), .B2(n17508), .ZN(
        n1339) );
  OAI221_X1 U1729 ( .B1(n18113), .B2(n18633), .C1(n19328), .C2(n18630), .A(
        n1329), .ZN(n1324) );
  AOI22_X1 U1730 ( .A1(n18627), .A2(n19696), .B1(n18624), .B2(n19448), .ZN(
        n1329) );
  OAI221_X1 U1731 ( .B1(n18081), .B2(n18681), .C1(n19312), .C2(n18678), .A(
        n1321), .ZN(n1316) );
  AOI22_X1 U1732 ( .A1(n18675), .A2(n19424), .B1(n18672), .B2(n17509), .ZN(
        n1321) );
  OAI221_X1 U1733 ( .B1(n18114), .B2(n18633), .C1(n19327), .C2(n18630), .A(
        n1311), .ZN(n1306) );
  AOI22_X1 U1734 ( .A1(n18627), .A2(n19695), .B1(n18624), .B2(n19447), .ZN(
        n1311) );
  OAI221_X1 U1735 ( .B1(n18082), .B2(n18681), .C1(n19311), .C2(n18678), .A(
        n1303), .ZN(n1298) );
  AOI22_X1 U1736 ( .A1(n18675), .A2(n19423), .B1(n18672), .B2(n17510), .ZN(
        n1303) );
  OAI221_X1 U1737 ( .B1(n18115), .B2(n18633), .C1(n18043), .C2(n18630), .A(
        n1293), .ZN(n1288) );
  AOI22_X1 U1738 ( .A1(n18627), .A2(n19694), .B1(n18624), .B2(n19446), .ZN(
        n1293) );
  OAI221_X1 U1739 ( .B1(n18083), .B2(n18681), .C1(n19310), .C2(n18678), .A(
        n1285), .ZN(n1280) );
  AOI22_X1 U1740 ( .A1(n18675), .A2(n19422), .B1(n18672), .B2(n17511), .ZN(
        n1285) );
  OAI221_X1 U1741 ( .B1(n18119), .B2(n18633), .C1(n18047), .C2(n18630), .A(
        n1221), .ZN(n1216) );
  AOI22_X1 U1742 ( .A1(n18627), .A2(n19690), .B1(n18623), .B2(n19442), .ZN(
        n1221) );
  OAI221_X1 U1743 ( .B1(n18087), .B2(n18681), .C1(n18063), .C2(n18678), .A(
        n1213), .ZN(n1208) );
  AOI22_X1 U1744 ( .A1(n18675), .A2(n19418), .B1(n18671), .B2(n17515), .ZN(
        n1213) );
  OAI221_X1 U1745 ( .B1(n18120), .B2(n18633), .C1(n19321), .C2(n18630), .A(
        n1203), .ZN(n1198) );
  AOI22_X1 U1746 ( .A1(n18627), .A2(n19689), .B1(n18623), .B2(n19441), .ZN(
        n1203) );
  OAI221_X1 U1747 ( .B1(n18088), .B2(n18681), .C1(n19305), .C2(n18678), .A(
        n1195), .ZN(n1190) );
  AOI22_X1 U1748 ( .A1(n18675), .A2(n19417), .B1(n18671), .B2(n17516), .ZN(
        n1195) );
  OAI221_X1 U1749 ( .B1(n18121), .B2(n18633), .C1(n19320), .C2(n18630), .A(
        n1185), .ZN(n1180) );
  AOI22_X1 U1750 ( .A1(n18627), .A2(n19688), .B1(n18623), .B2(n19440), .ZN(
        n1185) );
  OAI221_X1 U1751 ( .B1(n18089), .B2(n18681), .C1(n19304), .C2(n18678), .A(
        n1177), .ZN(n1172) );
  AOI22_X1 U1752 ( .A1(n18675), .A2(n19416), .B1(n18671), .B2(n17517), .ZN(
        n1177) );
  OAI221_X1 U1753 ( .B1(n18122), .B2(n18633), .C1(n19319), .C2(n18630), .A(
        n1167), .ZN(n1162) );
  AOI22_X1 U1754 ( .A1(n18627), .A2(n19687), .B1(n18623), .B2(n19439), .ZN(
        n1167) );
  OAI221_X1 U1755 ( .B1(n18090), .B2(n18681), .C1(n19303), .C2(n18678), .A(
        n1159), .ZN(n1154) );
  AOI22_X1 U1756 ( .A1(n18675), .A2(n19415), .B1(n18671), .B2(n17518), .ZN(
        n1159) );
  OAI221_X1 U1757 ( .B1(n18105), .B2(n18632), .C1(n19336), .C2(n18629), .A(
        n1473), .ZN(n1468) );
  AOI22_X1 U1758 ( .A1(n18626), .A2(n19608), .B1(n18625), .B2(n19456), .ZN(
        n1473) );
  OAI221_X1 U1759 ( .B1(n18289), .B2(n18680), .C1(n19200), .C2(n18677), .A(
        n1465), .ZN(n1460) );
  AOI22_X1 U1760 ( .A1(n18674), .A2(n19432), .B1(n18673), .B2(n17661), .ZN(
        n1465) );
  OAI221_X1 U1761 ( .B1(n18106), .B2(n18632), .C1(n19335), .C2(n18629), .A(
        n1455), .ZN(n1450) );
  AOI22_X1 U1762 ( .A1(n18626), .A2(n19607), .B1(n18625), .B2(n19455), .ZN(
        n1455) );
  OAI221_X1 U1763 ( .B1(n18290), .B2(n18680), .C1(n19199), .C2(n18677), .A(
        n1447), .ZN(n1442) );
  AOI22_X1 U1764 ( .A1(n18674), .A2(n19431), .B1(n18673), .B2(n17662), .ZN(
        n1447) );
  OAI221_X1 U1765 ( .B1(n18107), .B2(n18632), .C1(n19334), .C2(n18629), .A(
        n1437), .ZN(n1432) );
  AOI22_X1 U1766 ( .A1(n18626), .A2(n19702), .B1(n18624), .B2(n19454), .ZN(
        n1437) );
  OAI221_X1 U1767 ( .B1(n18075), .B2(n18680), .C1(n19318), .C2(n18677), .A(
        n1429), .ZN(n1424) );
  AOI22_X1 U1768 ( .A1(n18674), .A2(n19430), .B1(n18672), .B2(n17503), .ZN(
        n1429) );
  OAI221_X1 U1769 ( .B1(n18108), .B2(n18632), .C1(n19333), .C2(n18629), .A(
        n1419), .ZN(n1414) );
  AOI22_X1 U1770 ( .A1(n18626), .A2(n19701), .B1(n18624), .B2(n19453), .ZN(
        n1419) );
  OAI221_X1 U1771 ( .B1(n18076), .B2(n18680), .C1(n19317), .C2(n18677), .A(
        n1411), .ZN(n1406) );
  AOI22_X1 U1772 ( .A1(n18674), .A2(n19429), .B1(n18672), .B2(n17504), .ZN(
        n1411) );
  OAI221_X1 U1773 ( .B1(n18102), .B2(n18632), .C1(n19339), .C2(n18629), .A(
        n1527), .ZN(n1522) );
  AOI22_X1 U1774 ( .A1(n18626), .A2(n19611), .B1(n18625), .B2(n19459), .ZN(
        n1527) );
  OAI221_X1 U1775 ( .B1(n18286), .B2(n18680), .C1(n19203), .C2(n18677), .A(
        n1519), .ZN(n1514) );
  AOI22_X1 U1776 ( .A1(n18674), .A2(n19435), .B1(n18673), .B2(n17658), .ZN(
        n1519) );
  OAI221_X1 U1777 ( .B1(n18298), .B2(n18634), .C1(n19207), .C2(n18631), .A(
        n1017), .ZN(n1002) );
  AOI22_X1 U1778 ( .A1(n18628), .A2(n19679), .B1(n18623), .B2(n19247), .ZN(
        n1017) );
  OAI221_X1 U1779 ( .B1(n18098), .B2(n18682), .C1(n19295), .C2(n18679), .A(
        n993), .ZN(n978) );
  AOI22_X1 U1780 ( .A1(n18676), .A2(n19239), .B1(n18671), .B2(n17526), .ZN(
        n993) );
  OAI221_X1 U1781 ( .B1(n18103), .B2(n18632), .C1(n18031), .C2(n18629), .A(
        n1509), .ZN(n1504) );
  AOI22_X1 U1782 ( .A1(n18626), .A2(n19610), .B1(n18625), .B2(n19458), .ZN(
        n1509) );
  OAI221_X1 U1783 ( .B1(n18287), .B2(n18680), .C1(n19202), .C2(n18677), .A(
        n1501), .ZN(n1496) );
  AOI22_X1 U1784 ( .A1(n18674), .A2(n19434), .B1(n18673), .B2(n17659), .ZN(
        n1501) );
  OAI221_X1 U1785 ( .B1(n18104), .B2(n18632), .C1(n19337), .C2(n18629), .A(
        n1491), .ZN(n1486) );
  AOI22_X1 U1786 ( .A1(n18626), .A2(n19609), .B1(n18625), .B2(n19457), .ZN(
        n1491) );
  OAI221_X1 U1787 ( .B1(n18288), .B2(n18680), .C1(n19201), .C2(n18677), .A(
        n1483), .ZN(n1478) );
  AOI22_X1 U1788 ( .A1(n18674), .A2(n19433), .B1(n18673), .B2(n17660), .ZN(
        n1483) );
  OAI221_X1 U1789 ( .B1(n18295), .B2(n18634), .C1(n19210), .C2(n18631), .A(
        n1077), .ZN(n1072) );
  AOI22_X1 U1790 ( .A1(n18628), .A2(n19682), .B1(n18623), .B2(n19250), .ZN(
        n1077) );
  OAI221_X1 U1791 ( .B1(n18095), .B2(n18682), .C1(n19298), .C2(n18679), .A(
        n1069), .ZN(n1064) );
  AOI22_X1 U1792 ( .A1(n18676), .A2(n19242), .B1(n18671), .B2(n17523), .ZN(
        n1069) );
  OAI221_X1 U1793 ( .B1(n18296), .B2(n18634), .C1(n19209), .C2(n18631), .A(
        n1059), .ZN(n1054) );
  AOI22_X1 U1794 ( .A1(n18628), .A2(n19681), .B1(n18623), .B2(n19249), .ZN(
        n1059) );
  OAI221_X1 U1795 ( .B1(n18096), .B2(n18682), .C1(n19297), .C2(n18679), .A(
        n1051), .ZN(n1046) );
  AOI22_X1 U1796 ( .A1(n18676), .A2(n19241), .B1(n18671), .B2(n17524), .ZN(
        n1051) );
  OAI221_X1 U1797 ( .B1(n18101), .B2(n18632), .C1(n19340), .C2(n18629), .A(
        n1545), .ZN(n1540) );
  AOI22_X1 U1798 ( .A1(n18626), .A2(n19612), .B1(n18625), .B2(n19460), .ZN(
        n1545) );
  OAI221_X1 U1799 ( .B1(n18285), .B2(n18680), .C1(n19204), .C2(n18677), .A(
        n1537), .ZN(n1532) );
  AOI22_X1 U1800 ( .A1(n18674), .A2(n19436), .B1(n18673), .B2(n17657), .ZN(
        n1537) );
  OAI221_X1 U1801 ( .B1(n18297), .B2(n18634), .C1(n19208), .C2(n18631), .A(
        n1041), .ZN(n1036) );
  AOI22_X1 U1802 ( .A1(n18628), .A2(n19680), .B1(n18623), .B2(n19248), .ZN(
        n1041) );
  OAI221_X1 U1803 ( .B1(n18097), .B2(n18682), .C1(n19296), .C2(n18679), .A(
        n1033), .ZN(n1028) );
  AOI22_X1 U1804 ( .A1(n18676), .A2(n19240), .B1(n18671), .B2(n17525), .ZN(
        n1033) );
  OAI221_X1 U1805 ( .B1(n18291), .B2(n18634), .C1(n19214), .C2(n18631), .A(
        n1149), .ZN(n1144) );
  AOI22_X1 U1806 ( .A1(n18628), .A2(n19686), .B1(n18623), .B2(n19254), .ZN(
        n1149) );
  OAI221_X1 U1807 ( .B1(n18091), .B2(n18682), .C1(n19302), .C2(n18679), .A(
        n1141), .ZN(n1136) );
  AOI22_X1 U1808 ( .A1(n18676), .A2(n19246), .B1(n18671), .B2(n17519), .ZN(
        n1141) );
  OAI221_X1 U1809 ( .B1(n18292), .B2(n18634), .C1(n19213), .C2(n18631), .A(
        n1131), .ZN(n1126) );
  AOI22_X1 U1810 ( .A1(n18628), .A2(n19685), .B1(n18623), .B2(n19253), .ZN(
        n1131) );
  OAI221_X1 U1811 ( .B1(n18092), .B2(n18682), .C1(n19301), .C2(n18679), .A(
        n1123), .ZN(n1118) );
  AOI22_X1 U1812 ( .A1(n18676), .A2(n19245), .B1(n18671), .B2(n17520), .ZN(
        n1123) );
  OAI221_X1 U1813 ( .B1(n18293), .B2(n18634), .C1(n19212), .C2(n18631), .A(
        n1113), .ZN(n1108) );
  AOI22_X1 U1814 ( .A1(n18628), .A2(n19684), .B1(n18623), .B2(n19252), .ZN(
        n1113) );
  OAI221_X1 U1815 ( .B1(n18093), .B2(n18682), .C1(n19300), .C2(n18679), .A(
        n1105), .ZN(n1100) );
  AOI22_X1 U1816 ( .A1(n18676), .A2(n19244), .B1(n18671), .B2(n17521), .ZN(
        n1105) );
  OAI221_X1 U1817 ( .B1(n18294), .B2(n18634), .C1(n19211), .C2(n18631), .A(
        n1095), .ZN(n1090) );
  AOI22_X1 U1818 ( .A1(n18628), .A2(n19683), .B1(n18623), .B2(n19251), .ZN(
        n1095) );
  OAI221_X1 U1819 ( .B1(n18094), .B2(n18682), .C1(n19299), .C2(n18679), .A(
        n1087), .ZN(n1082) );
  AOI22_X1 U1820 ( .A1(n18676), .A2(n19243), .B1(n18671), .B2(n17522), .ZN(
        n1087) );
  OAI221_X1 U1821 ( .B1(n17855), .B2(n18536), .C1(n18131), .C2(n18533), .A(
        n2057), .ZN(n2052) );
  AOI22_X1 U1822 ( .A1(n18530), .A2(n18035), .B1(n18528), .B2(n19702), .ZN(
        n2057) );
  OAI221_X1 U1823 ( .B1(n17856), .B2(n18536), .C1(n18132), .C2(n18533), .A(
        n2039), .ZN(n2034) );
  AOI22_X1 U1824 ( .A1(n18530), .A2(n18036), .B1(n18528), .B2(n19701), .ZN(
        n2039) );
  OAI221_X1 U1825 ( .B1(n17857), .B2(n18536), .C1(n18133), .C2(n18533), .A(
        n2021), .ZN(n2016) );
  AOI22_X1 U1826 ( .A1(n18530), .A2(n18037), .B1(n18528), .B2(n19700), .ZN(
        n2021) );
  OAI221_X1 U1827 ( .B1(n17858), .B2(n18536), .C1(n18134), .C2(n18533), .A(
        n2003), .ZN(n1998) );
  AOI22_X1 U1828 ( .A1(n18530), .A2(n18038), .B1(n18528), .B2(n19699), .ZN(
        n2003) );
  OAI221_X1 U1829 ( .B1(n17859), .B2(n18537), .C1(n18135), .C2(n18534), .A(
        n1985), .ZN(n1980) );
  AOI22_X1 U1830 ( .A1(n18531), .A2(n18039), .B1(n18528), .B2(n19698), .ZN(
        n1985) );
  OAI221_X1 U1831 ( .B1(n17860), .B2(n18537), .C1(n18136), .C2(n18534), .A(
        n1967), .ZN(n1962) );
  AOI22_X1 U1832 ( .A1(n18531), .A2(n18040), .B1(n18528), .B2(n19697), .ZN(
        n1967) );
  OAI221_X1 U1833 ( .B1(n17861), .B2(n18537), .C1(n18137), .C2(n18534), .A(
        n1949), .ZN(n1944) );
  AOI22_X1 U1834 ( .A1(n18531), .A2(n18041), .B1(n18528), .B2(n19696), .ZN(
        n1949) );
  OAI221_X1 U1835 ( .B1(n17862), .B2(n18537), .C1(n18138), .C2(n18534), .A(
        n1931), .ZN(n1926) );
  AOI22_X1 U1836 ( .A1(n18531), .A2(n18042), .B1(n18528), .B2(n19695), .ZN(
        n1931) );
  OAI221_X1 U1837 ( .B1(n17863), .B2(n18537), .C1(n18139), .C2(n18534), .A(
        n1913), .ZN(n1908) );
  AOI22_X1 U1838 ( .A1(n18531), .A2(n19326), .B1(n18528), .B2(n19694), .ZN(
        n1913) );
  OAI221_X1 U1839 ( .B1(n17864), .B2(n18537), .C1(n18140), .C2(n18534), .A(
        n1895), .ZN(n1890) );
  AOI22_X1 U1840 ( .A1(n18531), .A2(n18044), .B1(n18528), .B2(n19693), .ZN(
        n1895) );
  OAI221_X1 U1841 ( .B1(n17865), .B2(n18537), .C1(n18141), .C2(n18534), .A(
        n1877), .ZN(n1872) );
  AOI22_X1 U1842 ( .A1(n18531), .A2(n19324), .B1(n18528), .B2(n19692), .ZN(
        n1877) );
  OAI221_X1 U1843 ( .B1(n17866), .B2(n18537), .C1(n18142), .C2(n18534), .A(
        n1859), .ZN(n1854) );
  AOI22_X1 U1844 ( .A1(n18531), .A2(n18046), .B1(n18528), .B2(n19691), .ZN(
        n1859) );
  OAI221_X1 U1845 ( .B1(n17867), .B2(n18537), .C1(n18143), .C2(n18534), .A(
        n1841), .ZN(n1836) );
  AOI22_X1 U1846 ( .A1(n18531), .A2(n19322), .B1(n18527), .B2(n19690), .ZN(
        n1841) );
  OAI221_X1 U1847 ( .B1(n17868), .B2(n18537), .C1(n18144), .C2(n18534), .A(
        n1823), .ZN(n1818) );
  AOI22_X1 U1848 ( .A1(n18531), .A2(n18048), .B1(n18527), .B2(n19689), .ZN(
        n1823) );
  OAI221_X1 U1849 ( .B1(n17869), .B2(n18537), .C1(n18145), .C2(n18534), .A(
        n1805), .ZN(n1800) );
  AOI22_X1 U1850 ( .A1(n18531), .A2(n18049), .B1(n18527), .B2(n19688), .ZN(
        n1805) );
  OAI221_X1 U1851 ( .B1(n17870), .B2(n18537), .C1(n18146), .C2(n18534), .A(
        n1787), .ZN(n1782) );
  AOI22_X1 U1852 ( .A1(n18531), .A2(n18050), .B1(n18527), .B2(n19687), .ZN(
        n1787) );
  OAI221_X1 U1853 ( .B1(n18211), .B2(n18538), .C1(n18299), .C2(n18535), .A(
        n1769), .ZN(n1764) );
  AOI22_X1 U1854 ( .A1(n18532), .A2(n18267), .B1(n18527), .B2(n19686), .ZN(
        n1769) );
  OAI221_X1 U1855 ( .B1(n18212), .B2(n18538), .C1(n18300), .C2(n18535), .A(
        n1751), .ZN(n1746) );
  AOI22_X1 U1856 ( .A1(n18532), .A2(n18268), .B1(n18527), .B2(n19685), .ZN(
        n1751) );
  OAI221_X1 U1857 ( .B1(n18213), .B2(n18538), .C1(n18301), .C2(n18535), .A(
        n1733), .ZN(n1728) );
  AOI22_X1 U1858 ( .A1(n18532), .A2(n18269), .B1(n18527), .B2(n19684), .ZN(
        n1733) );
  OAI221_X1 U1859 ( .B1(n18214), .B2(n18538), .C1(n18302), .C2(n18535), .A(
        n1715), .ZN(n1710) );
  AOI22_X1 U1860 ( .A1(n18532), .A2(n18270), .B1(n18527), .B2(n19683), .ZN(
        n1715) );
  OAI221_X1 U1861 ( .B1(n18215), .B2(n18538), .C1(n18303), .C2(n18535), .A(
        n1697), .ZN(n1692) );
  AOI22_X1 U1862 ( .A1(n18532), .A2(n18271), .B1(n18527), .B2(n19682), .ZN(
        n1697) );
  OAI221_X1 U1863 ( .B1(n18216), .B2(n18538), .C1(n18304), .C2(n18535), .A(
        n1679), .ZN(n1674) );
  AOI22_X1 U1864 ( .A1(n18532), .A2(n18272), .B1(n18527), .B2(n19681), .ZN(
        n1679) );
  OAI221_X1 U1865 ( .B1(n18217), .B2(n18538), .C1(n18305), .C2(n18535), .A(
        n1661), .ZN(n1656) );
  AOI22_X1 U1866 ( .A1(n18532), .A2(n18273), .B1(n18527), .B2(n19680), .ZN(
        n1661) );
  OAI221_X1 U1867 ( .B1(n18218), .B2(n18538), .C1(n18306), .C2(n18535), .A(
        n1637), .ZN(n1622) );
  AOI22_X1 U1868 ( .A1(n18532), .A2(n18274), .B1(n18527), .B2(n19679), .ZN(
        n1637) );
  OAI221_X1 U1869 ( .B1(n17895), .B2(n18584), .C1(n17815), .C2(n18581), .A(
        n2202), .ZN(n2188) );
  AOI22_X1 U1870 ( .A1(n18578), .A2(n19542), .B1(n18577), .B2(n17647), .ZN(
        n2202) );
  OAI221_X1 U1871 ( .B1(n17896), .B2(n18584), .C1(n17816), .C2(n18581), .A(
        n2175), .ZN(n2170) );
  AOI22_X1 U1872 ( .A1(n18578), .A2(n19541), .B1(n18577), .B2(n17648), .ZN(
        n2175) );
  OAI221_X1 U1873 ( .B1(n17897), .B2(n18584), .C1(n17817), .C2(n18581), .A(
        n2157), .ZN(n2152) );
  AOI22_X1 U1874 ( .A1(n18578), .A2(n19540), .B1(n18577), .B2(n17649), .ZN(
        n2157) );
  OAI221_X1 U1875 ( .B1(n17898), .B2(n18584), .C1(n17818), .C2(n18581), .A(
        n2139), .ZN(n2134) );
  AOI22_X1 U1876 ( .A1(n18578), .A2(n19539), .B1(n18577), .B2(n17650), .ZN(
        n2139) );
  OAI221_X1 U1877 ( .B1(n17899), .B2(n18584), .C1(n17819), .C2(n18581), .A(
        n2121), .ZN(n2116) );
  AOI22_X1 U1878 ( .A1(n18578), .A2(n19538), .B1(n18577), .B2(n17651), .ZN(
        n2121) );
  OAI221_X1 U1879 ( .B1(n17900), .B2(n18584), .C1(n17820), .C2(n18581), .A(
        n2103), .ZN(n2098) );
  AOI22_X1 U1880 ( .A1(n18578), .A2(n19537), .B1(n18577), .B2(n17652), .ZN(
        n2103) );
  OAI221_X1 U1881 ( .B1(n17901), .B2(n18584), .C1(n17821), .C2(n18581), .A(
        n2085), .ZN(n2080) );
  AOI22_X1 U1882 ( .A1(n18578), .A2(n19536), .B1(n18577), .B2(n17653), .ZN(
        n2085) );
  OAI221_X1 U1883 ( .B1(n17902), .B2(n18584), .C1(n17822), .C2(n18581), .A(
        n2067), .ZN(n2062) );
  AOI22_X1 U1884 ( .A1(n18578), .A2(n19535), .B1(n18577), .B2(n17654), .ZN(
        n2067) );
  OAI221_X1 U1885 ( .B1(n18107), .B2(n18524), .C1(n19824), .C2(n18521), .A(
        n2058), .ZN(n2051) );
  AOI22_X1 U1886 ( .A1(n18518), .A2(n18346), .B1(n18516), .B2(n19414), .ZN(
        n2058) );
  OAI221_X1 U1887 ( .B1(n18108), .B2(n18524), .C1(n19823), .C2(n18521), .A(
        n2040), .ZN(n2033) );
  AOI22_X1 U1888 ( .A1(n18518), .A2(n18347), .B1(n18516), .B2(n19413), .ZN(
        n2040) );
  OAI221_X1 U1889 ( .B1(n18109), .B2(n18524), .C1(n17966), .C2(n18521), .A(
        n2022), .ZN(n2015) );
  AOI22_X1 U1890 ( .A1(n18518), .A2(n18348), .B1(n18516), .B2(n19412), .ZN(
        n2022) );
  OAI221_X1 U1891 ( .B1(n18110), .B2(n18524), .C1(n17967), .C2(n18521), .A(
        n2004), .ZN(n1997) );
  AOI22_X1 U1892 ( .A1(n18518), .A2(n18349), .B1(n18516), .B2(n19411), .ZN(
        n2004) );
  OAI221_X1 U1893 ( .B1(n18111), .B2(n18525), .C1(n17968), .C2(n18522), .A(
        n1986), .ZN(n1979) );
  AOI22_X1 U1894 ( .A1(n18519), .A2(n18350), .B1(n18516), .B2(n19410), .ZN(
        n1986) );
  OAI221_X1 U1895 ( .B1(n18112), .B2(n18525), .C1(n17969), .C2(n18522), .A(
        n1968), .ZN(n1961) );
  AOI22_X1 U1896 ( .A1(n18519), .A2(n18351), .B1(n18516), .B2(n19409), .ZN(
        n1968) );
  OAI221_X1 U1897 ( .B1(n18113), .B2(n18525), .C1(n17970), .C2(n18522), .A(
        n1950), .ZN(n1943) );
  AOI22_X1 U1898 ( .A1(n18519), .A2(n18352), .B1(n18516), .B2(n19408), .ZN(
        n1950) );
  OAI221_X1 U1899 ( .B1(n18114), .B2(n18525), .C1(n17971), .C2(n18522), .A(
        n1932), .ZN(n1925) );
  AOI22_X1 U1900 ( .A1(n18519), .A2(n18353), .B1(n18516), .B2(n19407), .ZN(
        n1932) );
  OAI221_X1 U1901 ( .B1(n18115), .B2(n18525), .C1(n17972), .C2(n18522), .A(
        n1914), .ZN(n1907) );
  AOI22_X1 U1902 ( .A1(n18519), .A2(n18354), .B1(n18516), .B2(n19406), .ZN(
        n1914) );
  OAI221_X1 U1903 ( .B1(n18116), .B2(n18525), .C1(n17973), .C2(n18522), .A(
        n1896), .ZN(n1889) );
  AOI22_X1 U1904 ( .A1(n18519), .A2(n18355), .B1(n18516), .B2(n19405), .ZN(
        n1896) );
  OAI221_X1 U1905 ( .B1(n18117), .B2(n18525), .C1(n17974), .C2(n18522), .A(
        n1878), .ZN(n1871) );
  AOI22_X1 U1906 ( .A1(n18519), .A2(n18356), .B1(n18516), .B2(n19404), .ZN(
        n1878) );
  OAI221_X1 U1907 ( .B1(n18118), .B2(n18525), .C1(n17975), .C2(n18522), .A(
        n1860), .ZN(n1853) );
  AOI22_X1 U1908 ( .A1(n18519), .A2(n18357), .B1(n18516), .B2(n19403), .ZN(
        n1860) );
  OAI221_X1 U1909 ( .B1(n18119), .B2(n18525), .C1(n17976), .C2(n18522), .A(
        n1842), .ZN(n1835) );
  AOI22_X1 U1910 ( .A1(n18519), .A2(n18358), .B1(n18515), .B2(n19402), .ZN(
        n1842) );
  OAI221_X1 U1911 ( .B1(n18120), .B2(n18525), .C1(n17977), .C2(n18522), .A(
        n1824), .ZN(n1817) );
  AOI22_X1 U1912 ( .A1(n18519), .A2(n18359), .B1(n18515), .B2(n19401), .ZN(
        n1824) );
  OAI221_X1 U1913 ( .B1(n18121), .B2(n18525), .C1(n17978), .C2(n18522), .A(
        n1806), .ZN(n1799) );
  AOI22_X1 U1914 ( .A1(n18519), .A2(n18360), .B1(n18515), .B2(n19400), .ZN(
        n1806) );
  OAI221_X1 U1915 ( .B1(n18122), .B2(n18525), .C1(n17979), .C2(n18522), .A(
        n1788), .ZN(n1781) );
  AOI22_X1 U1916 ( .A1(n18519), .A2(n18361), .B1(n18515), .B2(n19399), .ZN(
        n1788) );
  OAI221_X1 U1917 ( .B1(n18291), .B2(n18526), .C1(n19662), .C2(n18523), .A(
        n1770), .ZN(n1763) );
  AOI22_X1 U1918 ( .A1(n18520), .A2(n18362), .B1(n18515), .B2(n19398), .ZN(
        n1770) );
  OAI221_X1 U1919 ( .B1(n18292), .B2(n18526), .C1(n19661), .C2(n18523), .A(
        n1752), .ZN(n1745) );
  AOI22_X1 U1920 ( .A1(n18520), .A2(n18363), .B1(n18515), .B2(n19397), .ZN(
        n1752) );
  OAI221_X1 U1921 ( .B1(n18293), .B2(n18526), .C1(n19660), .C2(n18523), .A(
        n1734), .ZN(n1727) );
  AOI22_X1 U1922 ( .A1(n18520), .A2(n18364), .B1(n18515), .B2(n19396), .ZN(
        n1734) );
  OAI221_X1 U1923 ( .B1(n18294), .B2(n18526), .C1(n19659), .C2(n18523), .A(
        n1716), .ZN(n1709) );
  AOI22_X1 U1924 ( .A1(n18520), .A2(n18365), .B1(n18515), .B2(n19395), .ZN(
        n1716) );
  OAI221_X1 U1925 ( .B1(n18295), .B2(n18526), .C1(n19658), .C2(n18523), .A(
        n1698), .ZN(n1691) );
  AOI22_X1 U1926 ( .A1(n18520), .A2(n18366), .B1(n18515), .B2(n19394), .ZN(
        n1698) );
  OAI221_X1 U1927 ( .B1(n18296), .B2(n18526), .C1(n19657), .C2(n18523), .A(
        n1680), .ZN(n1673) );
  AOI22_X1 U1928 ( .A1(n18520), .A2(n18367), .B1(n18515), .B2(n19393), .ZN(
        n1680) );
  OAI221_X1 U1929 ( .B1(n18297), .B2(n18526), .C1(n19656), .C2(n18523), .A(
        n1662), .ZN(n1655) );
  AOI22_X1 U1930 ( .A1(n18520), .A2(n18368), .B1(n18515), .B2(n19392), .ZN(
        n1662) );
  OAI221_X1 U1931 ( .B1(n18298), .B2(n18526), .C1(n19655), .C2(n18523), .A(
        n1642), .ZN(n1621) );
  AOI22_X1 U1932 ( .A1(n18520), .A2(n18369), .B1(n18515), .B2(n19391), .ZN(
        n1642) );
  OAI221_X1 U1933 ( .B1(n19143), .B2(n18622), .C1(n17965), .C2(n18619), .A(
        n1022), .ZN(n1001) );
  AOI22_X1 U1934 ( .A1(n18616), .A2(n19775), .B1(n18611), .B2(n19263), .ZN(
        n1022) );
  OAI221_X1 U1935 ( .B1(n19146), .B2(n18622), .C1(n17962), .C2(n18619), .A(
        n1078), .ZN(n1071) );
  AOI22_X1 U1936 ( .A1(n18616), .A2(n19778), .B1(n18611), .B2(n19266), .ZN(
        n1078) );
  OAI221_X1 U1937 ( .B1(n19145), .B2(n18622), .C1(n17963), .C2(n18619), .A(
        n1060), .ZN(n1053) );
  AOI22_X1 U1938 ( .A1(n18616), .A2(n19777), .B1(n18611), .B2(n19265), .ZN(
        n1060) );
  OAI221_X1 U1939 ( .B1(n19144), .B2(n18622), .C1(n17964), .C2(n18619), .A(
        n1042), .ZN(n1035) );
  AOI22_X1 U1940 ( .A1(n18616), .A2(n19776), .B1(n18611), .B2(n19264), .ZN(
        n1042) );
  OAI221_X1 U1941 ( .B1(n19150), .B2(n18622), .C1(n17958), .C2(n18619), .A(
        n1150), .ZN(n1143) );
  AOI22_X1 U1942 ( .A1(n18616), .A2(n19782), .B1(n18611), .B2(n19270), .ZN(
        n1150) );
  OAI221_X1 U1943 ( .B1(n19149), .B2(n18622), .C1(n17959), .C2(n18619), .A(
        n1132), .ZN(n1125) );
  AOI22_X1 U1944 ( .A1(n18616), .A2(n19781), .B1(n18611), .B2(n19269), .ZN(
        n1132) );
  OAI221_X1 U1945 ( .B1(n19148), .B2(n18622), .C1(n17960), .C2(n18619), .A(
        n1114), .ZN(n1107) );
  AOI22_X1 U1946 ( .A1(n18616), .A2(n19780), .B1(n18611), .B2(n19268), .ZN(
        n1114) );
  OAI221_X1 U1947 ( .B1(n19147), .B2(n18622), .C1(n17961), .C2(n18619), .A(
        n1096), .ZN(n1089) );
  AOI22_X1 U1948 ( .A1(n18616), .A2(n19779), .B1(n18611), .B2(n19267), .ZN(
        n1096) );
  OAI221_X1 U1949 ( .B1(n19134), .B2(n18620), .C1(n18243), .C2(n18617), .A(
        n1594), .ZN(n1587) );
  AOI22_X1 U1950 ( .A1(n18614), .A2(n19646), .B1(n18613), .B2(n19518), .ZN(
        n1594) );
  OAI221_X1 U1951 ( .B1(n19164), .B2(n18620), .C1(n17944), .C2(n18617), .A(
        n1402), .ZN(n1395) );
  AOI22_X1 U1952 ( .A1(n18614), .A2(n19796), .B1(n18612), .B2(n19508), .ZN(
        n1402) );
  OAI221_X1 U1953 ( .B1(n19163), .B2(n18620), .C1(n17945), .C2(n18617), .A(
        n1384), .ZN(n1377) );
  AOI22_X1 U1954 ( .A1(n18614), .A2(n19795), .B1(n18612), .B2(n19507), .ZN(
        n1384) );
  OAI221_X1 U1955 ( .B1(n19162), .B2(n18621), .C1(n17946), .C2(n18618), .A(
        n1366), .ZN(n1359) );
  AOI22_X1 U1956 ( .A1(n18615), .A2(n19794), .B1(n18612), .B2(n19506), .ZN(
        n1366) );
  OAI221_X1 U1957 ( .B1(n19157), .B2(n18621), .C1(n17951), .C2(n18618), .A(
        n1276), .ZN(n1269) );
  AOI22_X1 U1958 ( .A1(n18615), .A2(n19789), .B1(n18612), .B2(n19501), .ZN(
        n1276) );
  OAI221_X1 U1959 ( .B1(n19156), .B2(n18621), .C1(n17952), .C2(n18618), .A(
        n1258), .ZN(n1251) );
  AOI22_X1 U1960 ( .A1(n18615), .A2(n19788), .B1(n18612), .B2(n19500), .ZN(
        n1258) );
  OAI221_X1 U1961 ( .B1(n19155), .B2(n18621), .C1(n17953), .C2(n18618), .A(
        n1240), .ZN(n1233) );
  AOI22_X1 U1962 ( .A1(n18615), .A2(n19787), .B1(n18612), .B2(n19499), .ZN(
        n1240) );
  OAI221_X1 U1963 ( .B1(n19133), .B2(n18620), .C1(n18244), .C2(n18617), .A(
        n1564), .ZN(n1557) );
  AOI22_X1 U1964 ( .A1(n18614), .A2(n19645), .B1(n18613), .B2(n19517), .ZN(
        n1564) );
  OAI221_X1 U1965 ( .B1(n19161), .B2(n18621), .C1(n17947), .C2(n18618), .A(
        n1348), .ZN(n1341) );
  AOI22_X1 U1966 ( .A1(n18615), .A2(n19793), .B1(n18612), .B2(n19505), .ZN(
        n1348) );
  OAI221_X1 U1967 ( .B1(n19160), .B2(n18621), .C1(n17948), .C2(n18618), .A(
        n1330), .ZN(n1323) );
  AOI22_X1 U1968 ( .A1(n18615), .A2(n19792), .B1(n18612), .B2(n19504), .ZN(
        n1330) );
  OAI221_X1 U1969 ( .B1(n19159), .B2(n18621), .C1(n17949), .C2(n18618), .A(
        n1312), .ZN(n1305) );
  AOI22_X1 U1970 ( .A1(n18615), .A2(n19791), .B1(n18612), .B2(n19503), .ZN(
        n1312) );
  OAI221_X1 U1971 ( .B1(n19158), .B2(n18621), .C1(n17950), .C2(n18618), .A(
        n1294), .ZN(n1287) );
  AOI22_X1 U1972 ( .A1(n18615), .A2(n19790), .B1(n18612), .B2(n19502), .ZN(
        n1294) );
  OAI221_X1 U1973 ( .B1(n19154), .B2(n18621), .C1(n17954), .C2(n18618), .A(
        n1222), .ZN(n1215) );
  AOI22_X1 U1974 ( .A1(n18615), .A2(n19786), .B1(n18611), .B2(n19498), .ZN(
        n1222) );
  OAI221_X1 U1975 ( .B1(n19153), .B2(n18621), .C1(n17955), .C2(n18618), .A(
        n1204), .ZN(n1197) );
  AOI22_X1 U1976 ( .A1(n18615), .A2(n19785), .B1(n18611), .B2(n19497), .ZN(
        n1204) );
  OAI221_X1 U1977 ( .B1(n19152), .B2(n18621), .C1(n17956), .C2(n18618), .A(
        n1186), .ZN(n1179) );
  AOI22_X1 U1978 ( .A1(n18615), .A2(n19784), .B1(n18611), .B2(n19496), .ZN(
        n1186) );
  OAI221_X1 U1979 ( .B1(n19151), .B2(n18621), .C1(n17957), .C2(n18618), .A(
        n1168), .ZN(n1161) );
  AOI22_X1 U1980 ( .A1(n18615), .A2(n19783), .B1(n18611), .B2(n19495), .ZN(
        n1168) );
  OAI221_X1 U1981 ( .B1(n19128), .B2(n18620), .C1(n18249), .C2(n18617), .A(
        n1474), .ZN(n1467) );
  AOI22_X1 U1982 ( .A1(n18614), .A2(n19640), .B1(n18613), .B2(n19512), .ZN(
        n1474) );
  OAI221_X1 U1983 ( .B1(n19127), .B2(n18620), .C1(n18250), .C2(n18617), .A(
        n1456), .ZN(n1449) );
  AOI22_X1 U1984 ( .A1(n18614), .A2(n19639), .B1(n18613), .B2(n19511), .ZN(
        n1456) );
  OAI221_X1 U1985 ( .B1(n19166), .B2(n18620), .C1(n17942), .C2(n18617), .A(
        n1438), .ZN(n1431) );
  AOI22_X1 U1986 ( .A1(n18614), .A2(n19798), .B1(n18612), .B2(n19510), .ZN(
        n1438) );
  OAI221_X1 U1987 ( .B1(n19165), .B2(n18620), .C1(n17943), .C2(n18617), .A(
        n1420), .ZN(n1413) );
  AOI22_X1 U1988 ( .A1(n18614), .A2(n19797), .B1(n18612), .B2(n19509), .ZN(
        n1420) );
  OAI221_X1 U1989 ( .B1(n19131), .B2(n18620), .C1(n18246), .C2(n18617), .A(
        n1528), .ZN(n1521) );
  AOI22_X1 U1990 ( .A1(n18614), .A2(n19643), .B1(n18613), .B2(n19515), .ZN(
        n1528) );
  OAI221_X1 U1991 ( .B1(n19130), .B2(n18620), .C1(n18247), .C2(n18617), .A(
        n1510), .ZN(n1503) );
  AOI22_X1 U1992 ( .A1(n18614), .A2(n19642), .B1(n18613), .B2(n19514), .ZN(
        n1510) );
  OAI221_X1 U1993 ( .B1(n19129), .B2(n18620), .C1(n18248), .C2(n18617), .A(
        n1492), .ZN(n1485) );
  AOI22_X1 U1994 ( .A1(n18614), .A2(n19641), .B1(n18613), .B2(n19513), .ZN(
        n1492) );
  OAI221_X1 U1995 ( .B1(n19132), .B2(n18620), .C1(n18245), .C2(n18617), .A(
        n1546), .ZN(n1539) );
  AOI22_X1 U1996 ( .A1(n18614), .A2(n19644), .B1(n18613), .B2(n19516), .ZN(
        n1546) );
  AND3_X1 U1997 ( .A1(n19916), .A2(n19915), .A3(RD1), .ZN(n1586) );
  AND3_X1 U1998 ( .A1(ADD_RD2[4]), .A2(n19919), .A3(RD2), .ZN(n2203) );
  AND3_X1 U1999 ( .A1(RD2), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n2192) );
  AND3_X1 U2000 ( .A1(RD2), .A2(n19918), .A3(ADD_RD2[3]), .ZN(n2210) );
  AND3_X1 U2001 ( .A1(n19919), .A2(n19918), .A3(RD2), .ZN(n2213) );
  OAI22_X1 U2002 ( .A1(n19049), .A2(n18440), .B1(n2280), .B2(n19046), .ZN(
        n9198) );
  OAI22_X1 U2003 ( .A1(n19049), .A2(n18437), .B1(n2271), .B2(n19047), .ZN(
        n9199) );
  OAI22_X1 U2004 ( .A1(n19049), .A2(n18434), .B1(n2262), .B2(n19046), .ZN(
        n9200) );
  OAI22_X1 U2005 ( .A1(n19048), .A2(n18431), .B1(n2253), .B2(n19047), .ZN(
        n9201) );
  OAI22_X1 U2006 ( .A1(n19048), .A2(n18428), .B1(n2244), .B2(n19046), .ZN(
        n9202) );
  OAI22_X1 U2007 ( .A1(n19048), .A2(n18425), .B1(n2235), .B2(n19047), .ZN(
        n9203) );
  OAI22_X1 U2008 ( .A1(n19048), .A2(n18422), .B1(n2226), .B2(n19046), .ZN(
        n9204) );
  OAI22_X1 U2009 ( .A1(n19048), .A2(n18419), .B1(n2217), .B2(n19047), .ZN(
        n9205) );
  AOI22_X1 U2010 ( .A1(n18530), .A2(n18027), .B1(n18529), .B2(n19614), .ZN(
        n2212) );
  AOI22_X1 U2011 ( .A1(n18542), .A2(n17703), .B1(n18541), .B2(n19230), .ZN(
        n2211) );
  AOI22_X1 U2012 ( .A1(n18518), .A2(n18378), .B1(n18517), .B2(n19238), .ZN(
        n2214) );
  AOI22_X1 U2013 ( .A1(n18530), .A2(n18028), .B1(n18529), .B2(n19613), .ZN(
        n2183) );
  AOI22_X1 U2014 ( .A1(n18542), .A2(n17704), .B1(n18541), .B2(n19229), .ZN(
        n2182) );
  AOI22_X1 U2015 ( .A1(n18518), .A2(n18379), .B1(n18517), .B2(n19237), .ZN(
        n2184) );
  AOI22_X1 U2016 ( .A1(n18530), .A2(n18029), .B1(n18529), .B2(n19612), .ZN(
        n2165) );
  AOI22_X1 U2017 ( .A1(n18542), .A2(n17705), .B1(n18541), .B2(n19228), .ZN(
        n2164) );
  AOI22_X1 U2018 ( .A1(n18518), .A2(n18380), .B1(n18517), .B2(n19236), .ZN(
        n2166) );
  AOI22_X1 U2019 ( .A1(n18530), .A2(n18030), .B1(n18529), .B2(n19611), .ZN(
        n2147) );
  AOI22_X1 U2020 ( .A1(n18542), .A2(n17706), .B1(n18541), .B2(n19227), .ZN(
        n2146) );
  AOI22_X1 U2021 ( .A1(n18518), .A2(n18381), .B1(n18517), .B2(n19235), .ZN(
        n2148) );
  AOI22_X1 U2022 ( .A1(n18530), .A2(n19338), .B1(n18529), .B2(n19610), .ZN(
        n2129) );
  AOI22_X1 U2023 ( .A1(n18542), .A2(n17707), .B1(n18541), .B2(n19226), .ZN(
        n2128) );
  AOI22_X1 U2024 ( .A1(n18518), .A2(n18382), .B1(n18517), .B2(n19234), .ZN(
        n2130) );
  AOI22_X1 U2025 ( .A1(n18530), .A2(n18032), .B1(n18529), .B2(n19609), .ZN(
        n2111) );
  AOI22_X1 U2026 ( .A1(n18542), .A2(n17708), .B1(n18541), .B2(n19225), .ZN(
        n2110) );
  AOI22_X1 U2027 ( .A1(n18518), .A2(n18383), .B1(n18517), .B2(n19233), .ZN(
        n2112) );
  AOI22_X1 U2028 ( .A1(n18530), .A2(n18033), .B1(n18529), .B2(n19608), .ZN(
        n2093) );
  AOI22_X1 U2029 ( .A1(n18542), .A2(n17709), .B1(n18541), .B2(n19224), .ZN(
        n2092) );
  AOI22_X1 U2030 ( .A1(n18518), .A2(n18384), .B1(n18517), .B2(n19232), .ZN(
        n2094) );
  AOI22_X1 U2031 ( .A1(n18530), .A2(n18034), .B1(n18529), .B2(n19607), .ZN(
        n2075) );
  AOI22_X1 U2032 ( .A1(n18542), .A2(n17710), .B1(n18541), .B2(n19223), .ZN(
        n2074) );
  AOI22_X1 U2033 ( .A1(n18518), .A2(n18385), .B1(n18517), .B2(n19231), .ZN(
        n2076) );
  AOI22_X1 U2034 ( .A1(n18590), .A2(n17599), .B1(n18588), .B2(n19358), .ZN(
        n2048) );
  AOI22_X1 U2035 ( .A1(n18578), .A2(n19534), .B1(n18576), .B2(n17479), .ZN(
        n2049) );
  AOI22_X1 U2036 ( .A1(n18566), .A2(n19182), .B1(n18564), .B2(n19798), .ZN(
        n2050) );
  AOI22_X1 U2037 ( .A1(n18590), .A2(n17600), .B1(n18588), .B2(n19357), .ZN(
        n2030) );
  AOI22_X1 U2038 ( .A1(n18578), .A2(n19533), .B1(n18576), .B2(n17480), .ZN(
        n2031) );
  AOI22_X1 U2039 ( .A1(n18566), .A2(n19181), .B1(n18564), .B2(n19797), .ZN(
        n2032) );
  AOI22_X1 U2040 ( .A1(n18590), .A2(n17601), .B1(n18588), .B2(n19356), .ZN(
        n2012) );
  AOI22_X1 U2041 ( .A1(n18578), .A2(n19532), .B1(n18576), .B2(n17481), .ZN(
        n2013) );
  AOI22_X1 U2042 ( .A1(n18566), .A2(n19180), .B1(n18564), .B2(n19796), .ZN(
        n2014) );
  AOI22_X1 U2043 ( .A1(n18590), .A2(n17602), .B1(n18588), .B2(n19355), .ZN(
        n1994) );
  AOI22_X1 U2044 ( .A1(n18578), .A2(n19531), .B1(n18576), .B2(n17482), .ZN(
        n1995) );
  AOI22_X1 U2045 ( .A1(n18566), .A2(n19179), .B1(n18564), .B2(n19795), .ZN(
        n1996) );
  AOI22_X1 U2046 ( .A1(n18591), .A2(n17603), .B1(n18588), .B2(n19354), .ZN(
        n1976) );
  AOI22_X1 U2047 ( .A1(n18579), .A2(n19530), .B1(n18576), .B2(n17483), .ZN(
        n1977) );
  AOI22_X1 U2048 ( .A1(n18567), .A2(n19178), .B1(n18564), .B2(n19794), .ZN(
        n1978) );
  AOI22_X1 U2049 ( .A1(n18591), .A2(n17604), .B1(n18588), .B2(n19353), .ZN(
        n1958) );
  AOI22_X1 U2050 ( .A1(n18579), .A2(n19529), .B1(n18576), .B2(n17484), .ZN(
        n1959) );
  AOI22_X1 U2051 ( .A1(n18567), .A2(n19177), .B1(n18564), .B2(n19793), .ZN(
        n1960) );
  AOI22_X1 U2052 ( .A1(n18591), .A2(n17605), .B1(n18588), .B2(n19352), .ZN(
        n1940) );
  AOI22_X1 U2053 ( .A1(n18579), .A2(n19528), .B1(n18576), .B2(n17485), .ZN(
        n1941) );
  AOI22_X1 U2054 ( .A1(n18567), .A2(n19176), .B1(n18564), .B2(n19792), .ZN(
        n1942) );
  AOI22_X1 U2055 ( .A1(n18591), .A2(n17606), .B1(n18588), .B2(n19351), .ZN(
        n1922) );
  AOI22_X1 U2056 ( .A1(n18579), .A2(n19527), .B1(n18576), .B2(n17486), .ZN(
        n1923) );
  AOI22_X1 U2057 ( .A1(n18567), .A2(n19175), .B1(n18564), .B2(n19791), .ZN(
        n1924) );
  AOI22_X1 U2058 ( .A1(n18591), .A2(n17607), .B1(n18588), .B2(n19350), .ZN(
        n1904) );
  AOI22_X1 U2059 ( .A1(n18579), .A2(n19526), .B1(n18576), .B2(n17487), .ZN(
        n1905) );
  AOI22_X1 U2060 ( .A1(n18567), .A2(n19174), .B1(n18564), .B2(n19790), .ZN(
        n1906) );
  AOI22_X1 U2061 ( .A1(n18591), .A2(n17608), .B1(n18588), .B2(n19349), .ZN(
        n1886) );
  AOI22_X1 U2062 ( .A1(n18579), .A2(n19525), .B1(n18576), .B2(n17488), .ZN(
        n1887) );
  AOI22_X1 U2063 ( .A1(n18567), .A2(n19173), .B1(n18564), .B2(n19789), .ZN(
        n1888) );
  AOI22_X1 U2064 ( .A1(n18591), .A2(n17609), .B1(n18588), .B2(n19348), .ZN(
        n1868) );
  AOI22_X1 U2065 ( .A1(n18579), .A2(n19524), .B1(n18576), .B2(n17489), .ZN(
        n1869) );
  AOI22_X1 U2066 ( .A1(n18567), .A2(n19172), .B1(n18564), .B2(n19788), .ZN(
        n1870) );
  AOI22_X1 U2067 ( .A1(n18591), .A2(n17610), .B1(n18588), .B2(n19347), .ZN(
        n1850) );
  AOI22_X1 U2068 ( .A1(n18579), .A2(n19523), .B1(n18576), .B2(n17490), .ZN(
        n1851) );
  AOI22_X1 U2069 ( .A1(n18567), .A2(n19171), .B1(n18564), .B2(n19787), .ZN(
        n1852) );
  AOI22_X1 U2070 ( .A1(n18591), .A2(n17611), .B1(n18587), .B2(n19346), .ZN(
        n1832) );
  AOI22_X1 U2071 ( .A1(n18579), .A2(n19522), .B1(n18575), .B2(n17491), .ZN(
        n1833) );
  AOI22_X1 U2072 ( .A1(n18567), .A2(n19170), .B1(n18563), .B2(n19786), .ZN(
        n1834) );
  AOI22_X1 U2073 ( .A1(n18591), .A2(n17612), .B1(n18587), .B2(n19345), .ZN(
        n1814) );
  AOI22_X1 U2074 ( .A1(n18579), .A2(n19521), .B1(n18575), .B2(n17492), .ZN(
        n1815) );
  AOI22_X1 U2075 ( .A1(n18567), .A2(n19169), .B1(n18563), .B2(n19785), .ZN(
        n1816) );
  AOI22_X1 U2076 ( .A1(n18591), .A2(n17613), .B1(n18587), .B2(n19344), .ZN(
        n1796) );
  AOI22_X1 U2077 ( .A1(n18579), .A2(n19520), .B1(n18575), .B2(n17493), .ZN(
        n1797) );
  AOI22_X1 U2078 ( .A1(n18567), .A2(n19168), .B1(n18563), .B2(n19784), .ZN(
        n1798) );
  AOI22_X1 U2079 ( .A1(n18591), .A2(n17614), .B1(n18587), .B2(n19343), .ZN(
        n1778) );
  AOI22_X1 U2080 ( .A1(n18579), .A2(n19519), .B1(n18575), .B2(n17494), .ZN(
        n1779) );
  AOI22_X1 U2081 ( .A1(n18567), .A2(n19167), .B1(n18563), .B2(n19783), .ZN(
        n1780) );
  AOI22_X1 U2082 ( .A1(n18592), .A2(n17615), .B1(n18587), .B2(n19222), .ZN(
        n1760) );
  AOI22_X1 U2083 ( .A1(n18580), .A2(n19470), .B1(n18575), .B2(n17495), .ZN(
        n1761) );
  AOI22_X1 U2084 ( .A1(n18568), .A2(n19142), .B1(n18563), .B2(n19782), .ZN(
        n1762) );
  AOI22_X1 U2085 ( .A1(n18592), .A2(n17616), .B1(n18587), .B2(n19221), .ZN(
        n1742) );
  AOI22_X1 U2086 ( .A1(n18580), .A2(n19469), .B1(n18575), .B2(n17496), .ZN(
        n1743) );
  AOI22_X1 U2087 ( .A1(n18568), .A2(n19141), .B1(n18563), .B2(n19781), .ZN(
        n1744) );
  AOI22_X1 U2088 ( .A1(n18592), .A2(n17617), .B1(n18587), .B2(n19220), .ZN(
        n1724) );
  AOI22_X1 U2089 ( .A1(n18580), .A2(n19468), .B1(n18575), .B2(n17497), .ZN(
        n1725) );
  AOI22_X1 U2090 ( .A1(n18568), .A2(n19140), .B1(n18563), .B2(n19780), .ZN(
        n1726) );
  AOI22_X1 U2091 ( .A1(n18592), .A2(n17618), .B1(n18587), .B2(n19219), .ZN(
        n1706) );
  AOI22_X1 U2092 ( .A1(n18580), .A2(n19467), .B1(n18575), .B2(n17498), .ZN(
        n1707) );
  AOI22_X1 U2093 ( .A1(n18568), .A2(n19139), .B1(n18563), .B2(n19779), .ZN(
        n1708) );
  AOI22_X1 U2094 ( .A1(n18592), .A2(n17619), .B1(n18587), .B2(n19218), .ZN(
        n1688) );
  AOI22_X1 U2095 ( .A1(n18580), .A2(n19466), .B1(n18575), .B2(n17499), .ZN(
        n1689) );
  AOI22_X1 U2096 ( .A1(n18568), .A2(n19138), .B1(n18563), .B2(n19778), .ZN(
        n1690) );
  AOI22_X1 U2097 ( .A1(n18592), .A2(n17620), .B1(n18587), .B2(n19217), .ZN(
        n1670) );
  AOI22_X1 U2098 ( .A1(n18580), .A2(n19465), .B1(n18575), .B2(n17500), .ZN(
        n1671) );
  AOI22_X1 U2099 ( .A1(n18568), .A2(n19137), .B1(n18563), .B2(n19777), .ZN(
        n1672) );
  AOI22_X1 U2100 ( .A1(n18592), .A2(n17621), .B1(n18587), .B2(n19216), .ZN(
        n1652) );
  AOI22_X1 U2101 ( .A1(n18580), .A2(n19464), .B1(n18575), .B2(n17501), .ZN(
        n1653) );
  AOI22_X1 U2102 ( .A1(n18568), .A2(n19136), .B1(n18563), .B2(n19776), .ZN(
        n1654) );
  AOI22_X1 U2103 ( .A1(n18592), .A2(n17622), .B1(n18587), .B2(n19215), .ZN(
        n1608) );
  AOI22_X1 U2104 ( .A1(n18580), .A2(n19463), .B1(n18575), .B2(n17502), .ZN(
        n1613) );
  AOI22_X1 U2105 ( .A1(n18568), .A2(n19135), .B1(n18563), .B2(n19775), .ZN(
        n1618) );
  OAI221_X1 U2106 ( .B1(n18283), .B2(n18608), .C1(n19670), .C2(n18605), .A(
        n2191), .ZN(n2190) );
  AOI22_X1 U2107 ( .A1(n18602), .A2(n19438), .B1(n18601), .B2(n19888), .ZN(
        n2191) );
  OAI221_X1 U2108 ( .B1(n19550), .B2(n18596), .C1(n19630), .C2(n18593), .A(
        n2197), .ZN(n2189) );
  AOI22_X1 U2109 ( .A1(n18590), .A2(n17687), .B1(n18589), .B2(n19366), .ZN(
        n2197) );
  OAI221_X1 U2110 ( .B1(n17791), .B2(n18572), .C1(n19774), .C2(n18569), .A(
        n2204), .ZN(n2187) );
  AOI22_X1 U2111 ( .A1(n18566), .A2(n19190), .B1(n18565), .B2(n19646), .ZN(
        n2204) );
  OAI221_X1 U2112 ( .B1(n18284), .B2(n18608), .C1(n19669), .C2(n18605), .A(
        n2173), .ZN(n2172) );
  AOI22_X1 U2113 ( .A1(n18602), .A2(n19437), .B1(n18601), .B2(n19887), .ZN(
        n2173) );
  OAI221_X1 U2114 ( .B1(n19549), .B2(n18596), .C1(n19629), .C2(n18593), .A(
        n2174), .ZN(n2171) );
  AOI22_X1 U2115 ( .A1(n18590), .A2(n17688), .B1(n18589), .B2(n19365), .ZN(
        n2174) );
  OAI221_X1 U2116 ( .B1(n17792), .B2(n18572), .C1(n19773), .C2(n18569), .A(
        n2176), .ZN(n2169) );
  AOI22_X1 U2117 ( .A1(n18566), .A2(n19189), .B1(n18565), .B2(n19645), .ZN(
        n2176) );
  OAI221_X1 U2118 ( .B1(n18285), .B2(n18608), .C1(n19668), .C2(n18605), .A(
        n2155), .ZN(n2154) );
  AOI22_X1 U2119 ( .A1(n18602), .A2(n19436), .B1(n18601), .B2(n19886), .ZN(
        n2155) );
  OAI221_X1 U2120 ( .B1(n19548), .B2(n18596), .C1(n19628), .C2(n18593), .A(
        n2156), .ZN(n2153) );
  AOI22_X1 U2121 ( .A1(n18590), .A2(n17689), .B1(n18589), .B2(n19364), .ZN(
        n2156) );
  OAI221_X1 U2122 ( .B1(n17793), .B2(n18572), .C1(n19772), .C2(n18569), .A(
        n2158), .ZN(n2151) );
  AOI22_X1 U2123 ( .A1(n18566), .A2(n19188), .B1(n18565), .B2(n19644), .ZN(
        n2158) );
  OAI221_X1 U2124 ( .B1(n18286), .B2(n18608), .C1(n19667), .C2(n18605), .A(
        n2137), .ZN(n2136) );
  AOI22_X1 U2125 ( .A1(n18602), .A2(n19435), .B1(n18601), .B2(n19885), .ZN(
        n2137) );
  OAI221_X1 U2126 ( .B1(n19547), .B2(n18596), .C1(n19627), .C2(n18593), .A(
        n2138), .ZN(n2135) );
  AOI22_X1 U2127 ( .A1(n18590), .A2(n17690), .B1(n18589), .B2(n19363), .ZN(
        n2138) );
  OAI221_X1 U2128 ( .B1(n17794), .B2(n18572), .C1(n19771), .C2(n18569), .A(
        n2140), .ZN(n2133) );
  AOI22_X1 U2129 ( .A1(n18566), .A2(n19187), .B1(n18565), .B2(n19643), .ZN(
        n2140) );
  OAI221_X1 U2130 ( .B1(n18287), .B2(n18608), .C1(n19666), .C2(n18605), .A(
        n2119), .ZN(n2118) );
  AOI22_X1 U2131 ( .A1(n18602), .A2(n19434), .B1(n18601), .B2(n19884), .ZN(
        n2119) );
  OAI221_X1 U2132 ( .B1(n19546), .B2(n18596), .C1(n19626), .C2(n18593), .A(
        n2120), .ZN(n2117) );
  AOI22_X1 U2133 ( .A1(n18590), .A2(n17691), .B1(n18589), .B2(n19362), .ZN(
        n2120) );
  OAI221_X1 U2134 ( .B1(n17795), .B2(n18572), .C1(n19770), .C2(n18569), .A(
        n2122), .ZN(n2115) );
  AOI22_X1 U2135 ( .A1(n18566), .A2(n19186), .B1(n18565), .B2(n19642), .ZN(
        n2122) );
  OAI221_X1 U2136 ( .B1(n18288), .B2(n18608), .C1(n19665), .C2(n18605), .A(
        n2101), .ZN(n2100) );
  AOI22_X1 U2137 ( .A1(n18602), .A2(n19433), .B1(n18601), .B2(n19883), .ZN(
        n2101) );
  OAI221_X1 U2138 ( .B1(n19545), .B2(n18596), .C1(n19625), .C2(n18593), .A(
        n2102), .ZN(n2099) );
  AOI22_X1 U2139 ( .A1(n18590), .A2(n17692), .B1(n18589), .B2(n19361), .ZN(
        n2102) );
  OAI221_X1 U2140 ( .B1(n17796), .B2(n18572), .C1(n19769), .C2(n18569), .A(
        n2104), .ZN(n2097) );
  AOI22_X1 U2141 ( .A1(n18566), .A2(n19185), .B1(n18565), .B2(n19641), .ZN(
        n2104) );
  OAI221_X1 U2142 ( .B1(n18289), .B2(n18608), .C1(n19664), .C2(n18605), .A(
        n2083), .ZN(n2082) );
  AOI22_X1 U2143 ( .A1(n18602), .A2(n19432), .B1(n18601), .B2(n19882), .ZN(
        n2083) );
  OAI221_X1 U2144 ( .B1(n19544), .B2(n18596), .C1(n19624), .C2(n18593), .A(
        n2084), .ZN(n2081) );
  AOI22_X1 U2145 ( .A1(n18590), .A2(n17693), .B1(n18589), .B2(n19360), .ZN(
        n2084) );
  OAI221_X1 U2146 ( .B1(n17797), .B2(n18572), .C1(n19768), .C2(n18569), .A(
        n2086), .ZN(n2079) );
  AOI22_X1 U2147 ( .A1(n18566), .A2(n19184), .B1(n18565), .B2(n19640), .ZN(
        n2086) );
  OAI221_X1 U2148 ( .B1(n18290), .B2(n18608), .C1(n19663), .C2(n18605), .A(
        n2065), .ZN(n2064) );
  AOI22_X1 U2149 ( .A1(n18602), .A2(n19431), .B1(n18601), .B2(n19881), .ZN(
        n2065) );
  OAI221_X1 U2150 ( .B1(n19543), .B2(n18596), .C1(n19623), .C2(n18593), .A(
        n2066), .ZN(n2063) );
  AOI22_X1 U2151 ( .A1(n18590), .A2(n17694), .B1(n18589), .B2(n19359), .ZN(
        n2066) );
  OAI221_X1 U2152 ( .B1(n17798), .B2(n18572), .C1(n19767), .C2(n18569), .A(
        n2068), .ZN(n2061) );
  AOI22_X1 U2153 ( .A1(n18566), .A2(n19183), .B1(n18565), .B2(n19639), .ZN(
        n2068) );
  OAI221_X1 U2154 ( .B1(n18075), .B2(n18608), .C1(n19856), .C2(n18605), .A(
        n2047), .ZN(n2046) );
  AOI22_X1 U2155 ( .A1(n18602), .A2(n19430), .B1(n18600), .B2(n19912), .ZN(
        n2047) );
  OAI221_X1 U2156 ( .B1(n17879), .B2(n18560), .C1(n18179), .C2(n18557), .A(
        n2055), .ZN(n2054) );
  AOI22_X1 U2157 ( .A1(n18554), .A2(n18051), .B1(n18552), .B2(n19286), .ZN(
        n2055) );
  OAI221_X1 U2158 ( .B1(n19718), .B2(n18548), .C1(n19814), .C2(n18545), .A(
        n2056), .ZN(n2053) );
  AOI22_X1 U2159 ( .A1(n18542), .A2(n17711), .B1(n18540), .B2(n19390), .ZN(
        n2056) );
  OAI221_X1 U2160 ( .B1(n18076), .B2(n18608), .C1(n19855), .C2(n18605), .A(
        n2029), .ZN(n2028) );
  AOI22_X1 U2161 ( .A1(n18602), .A2(n19429), .B1(n18600), .B2(n19911), .ZN(
        n2029) );
  OAI221_X1 U2162 ( .B1(n17880), .B2(n18560), .C1(n18180), .C2(n18557), .A(
        n2037), .ZN(n2036) );
  AOI22_X1 U2163 ( .A1(n18554), .A2(n18052), .B1(n18552), .B2(n19285), .ZN(
        n2037) );
  OAI221_X1 U2164 ( .B1(n19717), .B2(n18548), .C1(n19813), .C2(n18545), .A(
        n2038), .ZN(n2035) );
  AOI22_X1 U2165 ( .A1(n18542), .A2(n17712), .B1(n18540), .B2(n19389), .ZN(
        n2038) );
  OAI221_X1 U2166 ( .B1(n18077), .B2(n18608), .C1(n19854), .C2(n18605), .A(
        n2011), .ZN(n2010) );
  AOI22_X1 U2167 ( .A1(n18602), .A2(n19428), .B1(n18600), .B2(n19910), .ZN(
        n2011) );
  OAI221_X1 U2168 ( .B1(n17881), .B2(n18560), .C1(n18181), .C2(n18557), .A(
        n2019), .ZN(n2018) );
  AOI22_X1 U2169 ( .A1(n18554), .A2(n18053), .B1(n18552), .B2(n19284), .ZN(
        n2019) );
  OAI221_X1 U2170 ( .B1(n19716), .B2(n18548), .C1(n19812), .C2(n18545), .A(
        n2020), .ZN(n2017) );
  AOI22_X1 U2171 ( .A1(n18542), .A2(n17713), .B1(n18540), .B2(n19388), .ZN(
        n2020) );
  OAI221_X1 U2172 ( .B1(n18078), .B2(n18608), .C1(n19853), .C2(n18605), .A(
        n1993), .ZN(n1992) );
  AOI22_X1 U2173 ( .A1(n18602), .A2(n19427), .B1(n18600), .B2(n19909), .ZN(
        n1993) );
  OAI221_X1 U2174 ( .B1(n17882), .B2(n18560), .C1(n18182), .C2(n18557), .A(
        n2001), .ZN(n2000) );
  AOI22_X1 U2175 ( .A1(n18554), .A2(n18054), .B1(n18552), .B2(n19283), .ZN(
        n2001) );
  OAI221_X1 U2176 ( .B1(n19715), .B2(n18548), .C1(n19811), .C2(n18545), .A(
        n2002), .ZN(n1999) );
  AOI22_X1 U2177 ( .A1(n18542), .A2(n17714), .B1(n18540), .B2(n19387), .ZN(
        n2002) );
  OAI221_X1 U2178 ( .B1(n18079), .B2(n18609), .C1(n19852), .C2(n18606), .A(
        n1975), .ZN(n1974) );
  AOI22_X1 U2179 ( .A1(n18603), .A2(n19426), .B1(n18600), .B2(n19908), .ZN(
        n1975) );
  OAI221_X1 U2180 ( .B1(n17883), .B2(n18561), .C1(n18183), .C2(n18558), .A(
        n1983), .ZN(n1982) );
  AOI22_X1 U2181 ( .A1(n18555), .A2(n18055), .B1(n18552), .B2(n19282), .ZN(
        n1983) );
  OAI221_X1 U2182 ( .B1(n19714), .B2(n18549), .C1(n19810), .C2(n18546), .A(
        n1984), .ZN(n1981) );
  AOI22_X1 U2183 ( .A1(n18543), .A2(n17715), .B1(n18540), .B2(n19386), .ZN(
        n1984) );
  OAI221_X1 U2184 ( .B1(n18080), .B2(n18609), .C1(n19851), .C2(n18606), .A(
        n1957), .ZN(n1956) );
  AOI22_X1 U2185 ( .A1(n18603), .A2(n19425), .B1(n18600), .B2(n19907), .ZN(
        n1957) );
  OAI221_X1 U2186 ( .B1(n17884), .B2(n18561), .C1(n18184), .C2(n18558), .A(
        n1965), .ZN(n1964) );
  AOI22_X1 U2187 ( .A1(n18555), .A2(n18056), .B1(n18552), .B2(n19281), .ZN(
        n1965) );
  OAI221_X1 U2188 ( .B1(n19713), .B2(n18549), .C1(n19809), .C2(n18546), .A(
        n1966), .ZN(n1963) );
  AOI22_X1 U2189 ( .A1(n18543), .A2(n17716), .B1(n18540), .B2(n19385), .ZN(
        n1966) );
  OAI221_X1 U2190 ( .B1(n18081), .B2(n18609), .C1(n19850), .C2(n18606), .A(
        n1939), .ZN(n1938) );
  AOI22_X1 U2191 ( .A1(n18603), .A2(n19424), .B1(n18600), .B2(n19906), .ZN(
        n1939) );
  OAI221_X1 U2192 ( .B1(n17885), .B2(n18561), .C1(n18185), .C2(n18558), .A(
        n1947), .ZN(n1946) );
  AOI22_X1 U2193 ( .A1(n18555), .A2(n18057), .B1(n18552), .B2(n19280), .ZN(
        n1947) );
  OAI221_X1 U2194 ( .B1(n19712), .B2(n18549), .C1(n19808), .C2(n18546), .A(
        n1948), .ZN(n1945) );
  AOI22_X1 U2195 ( .A1(n18543), .A2(n17717), .B1(n18540), .B2(n19384), .ZN(
        n1948) );
  OAI221_X1 U2196 ( .B1(n18082), .B2(n18609), .C1(n19849), .C2(n18606), .A(
        n1921), .ZN(n1920) );
  AOI22_X1 U2197 ( .A1(n18603), .A2(n19423), .B1(n18600), .B2(n19905), .ZN(
        n1921) );
  OAI221_X1 U2198 ( .B1(n17886), .B2(n18561), .C1(n18186), .C2(n18558), .A(
        n1929), .ZN(n1928) );
  AOI22_X1 U2199 ( .A1(n18555), .A2(n18058), .B1(n18552), .B2(n19279), .ZN(
        n1929) );
  OAI221_X1 U2200 ( .B1(n19711), .B2(n18549), .C1(n19807), .C2(n18546), .A(
        n1930), .ZN(n1927) );
  AOI22_X1 U2201 ( .A1(n18543), .A2(n17718), .B1(n18540), .B2(n19383), .ZN(
        n1930) );
  OAI221_X1 U2202 ( .B1(n18083), .B2(n18609), .C1(n19848), .C2(n18606), .A(
        n1903), .ZN(n1902) );
  AOI22_X1 U2203 ( .A1(n18603), .A2(n19422), .B1(n18600), .B2(n19904), .ZN(
        n1903) );
  OAI221_X1 U2204 ( .B1(n17887), .B2(n18561), .C1(n18187), .C2(n18558), .A(
        n1911), .ZN(n1910) );
  AOI22_X1 U2205 ( .A1(n18555), .A2(n18059), .B1(n18552), .B2(n19278), .ZN(
        n1911) );
  OAI221_X1 U2206 ( .B1(n19710), .B2(n18549), .C1(n19806), .C2(n18546), .A(
        n1912), .ZN(n1909) );
  AOI22_X1 U2207 ( .A1(n18543), .A2(n17719), .B1(n18540), .B2(n19382), .ZN(
        n1912) );
  OAI221_X1 U2208 ( .B1(n18084), .B2(n18609), .C1(n19847), .C2(n18606), .A(
        n1885), .ZN(n1884) );
  AOI22_X1 U2209 ( .A1(n18603), .A2(n19421), .B1(n18600), .B2(n19903), .ZN(
        n1885) );
  OAI221_X1 U2210 ( .B1(n17888), .B2(n18561), .C1(n18188), .C2(n18558), .A(
        n1893), .ZN(n1892) );
  AOI22_X1 U2211 ( .A1(n18555), .A2(n18060), .B1(n18552), .B2(n19277), .ZN(
        n1893) );
  OAI221_X1 U2212 ( .B1(n19709), .B2(n18549), .C1(n19805), .C2(n18546), .A(
        n1894), .ZN(n1891) );
  AOI22_X1 U2213 ( .A1(n18543), .A2(n17720), .B1(n18540), .B2(n19381), .ZN(
        n1894) );
  OAI221_X1 U2214 ( .B1(n18085), .B2(n18609), .C1(n19846), .C2(n18606), .A(
        n1867), .ZN(n1866) );
  AOI22_X1 U2215 ( .A1(n18603), .A2(n19420), .B1(n18600), .B2(n19902), .ZN(
        n1867) );
  OAI221_X1 U2216 ( .B1(n17889), .B2(n18561), .C1(n18189), .C2(n18558), .A(
        n1875), .ZN(n1874) );
  AOI22_X1 U2217 ( .A1(n18555), .A2(n18061), .B1(n18552), .B2(n19276), .ZN(
        n1875) );
  OAI221_X1 U2218 ( .B1(n19708), .B2(n18549), .C1(n19804), .C2(n18546), .A(
        n1876), .ZN(n1873) );
  AOI22_X1 U2219 ( .A1(n18543), .A2(n17721), .B1(n18540), .B2(n19380), .ZN(
        n1876) );
  OAI221_X1 U2220 ( .B1(n18086), .B2(n18609), .C1(n19845), .C2(n18606), .A(
        n1849), .ZN(n1848) );
  AOI22_X1 U2221 ( .A1(n18603), .A2(n19419), .B1(n18600), .B2(n19901), .ZN(
        n1849) );
  OAI221_X1 U2222 ( .B1(n17890), .B2(n18561), .C1(n18190), .C2(n18558), .A(
        n1857), .ZN(n1856) );
  AOI22_X1 U2223 ( .A1(n18555), .A2(n18062), .B1(n18552), .B2(n19275), .ZN(
        n1857) );
  OAI221_X1 U2224 ( .B1(n19707), .B2(n18549), .C1(n19803), .C2(n18546), .A(
        n1858), .ZN(n1855) );
  AOI22_X1 U2225 ( .A1(n18543), .A2(n17722), .B1(n18540), .B2(n19379), .ZN(
        n1858) );
  OAI221_X1 U2226 ( .B1(n18087), .B2(n18609), .C1(n19844), .C2(n18606), .A(
        n1831), .ZN(n1830) );
  AOI22_X1 U2227 ( .A1(n18603), .A2(n19418), .B1(n18599), .B2(n19900), .ZN(
        n1831) );
  OAI221_X1 U2228 ( .B1(n17891), .B2(n18561), .C1(n18191), .C2(n18558), .A(
        n1839), .ZN(n1838) );
  AOI22_X1 U2229 ( .A1(n18555), .A2(n19306), .B1(n18551), .B2(n19274), .ZN(
        n1839) );
  OAI221_X1 U2230 ( .B1(n19706), .B2(n18549), .C1(n19802), .C2(n18546), .A(
        n1840), .ZN(n1837) );
  AOI22_X1 U2231 ( .A1(n18543), .A2(n17723), .B1(n18539), .B2(n19378), .ZN(
        n1840) );
  OAI221_X1 U2232 ( .B1(n18088), .B2(n18609), .C1(n19843), .C2(n18606), .A(
        n1813), .ZN(n1812) );
  AOI22_X1 U2233 ( .A1(n18603), .A2(n19417), .B1(n18599), .B2(n19899), .ZN(
        n1813) );
  OAI221_X1 U2234 ( .B1(n17892), .B2(n18561), .C1(n18192), .C2(n18558), .A(
        n1821), .ZN(n1820) );
  AOI22_X1 U2235 ( .A1(n18555), .A2(n18064), .B1(n18551), .B2(n19273), .ZN(
        n1821) );
  OAI221_X1 U2236 ( .B1(n19705), .B2(n18549), .C1(n19801), .C2(n18546), .A(
        n1822), .ZN(n1819) );
  AOI22_X1 U2237 ( .A1(n18543), .A2(n17724), .B1(n18539), .B2(n19377), .ZN(
        n1822) );
  OAI221_X1 U2238 ( .B1(n18089), .B2(n18609), .C1(n19842), .C2(n18606), .A(
        n1795), .ZN(n1794) );
  AOI22_X1 U2239 ( .A1(n18603), .A2(n19416), .B1(n18599), .B2(n19898), .ZN(
        n1795) );
  OAI221_X1 U2240 ( .B1(n17893), .B2(n18561), .C1(n18193), .C2(n18558), .A(
        n1803), .ZN(n1802) );
  AOI22_X1 U2241 ( .A1(n18555), .A2(n18065), .B1(n18551), .B2(n19272), .ZN(
        n1803) );
  OAI221_X1 U2242 ( .B1(n19704), .B2(n18549), .C1(n19800), .C2(n18546), .A(
        n1804), .ZN(n1801) );
  AOI22_X1 U2243 ( .A1(n18543), .A2(n17725), .B1(n18539), .B2(n19376), .ZN(
        n1804) );
  OAI221_X1 U2244 ( .B1(n18090), .B2(n18609), .C1(n19841), .C2(n18606), .A(
        n1777), .ZN(n1776) );
  AOI22_X1 U2245 ( .A1(n18603), .A2(n19415), .B1(n18599), .B2(n19897), .ZN(
        n1777) );
  OAI221_X1 U2246 ( .B1(n17894), .B2(n18561), .C1(n18194), .C2(n18558), .A(
        n1785), .ZN(n1784) );
  AOI22_X1 U2247 ( .A1(n18555), .A2(n18066), .B1(n18551), .B2(n19271), .ZN(
        n1785) );
  OAI221_X1 U2248 ( .B1(n19703), .B2(n18549), .C1(n19799), .C2(n18546), .A(
        n1786), .ZN(n1783) );
  AOI22_X1 U2249 ( .A1(n18543), .A2(n17726), .B1(n18539), .B2(n19375), .ZN(
        n1786) );
  OAI221_X1 U2250 ( .B1(n19622), .B2(n18550), .C1(n19654), .C2(n18547), .A(
        n1768), .ZN(n1765) );
  AOI22_X1 U2251 ( .A1(n18544), .A2(n17751), .B1(n18539), .B2(n19374), .ZN(
        n1768) );
  OAI221_X1 U2252 ( .B1(n19621), .B2(n18550), .C1(n19653), .C2(n18547), .A(
        n1750), .ZN(n1747) );
  AOI22_X1 U2253 ( .A1(n18544), .A2(n17752), .B1(n18539), .B2(n19373), .ZN(
        n1750) );
  OAI221_X1 U2254 ( .B1(n19620), .B2(n18550), .C1(n19652), .C2(n18547), .A(
        n1732), .ZN(n1729) );
  AOI22_X1 U2255 ( .A1(n18544), .A2(n17753), .B1(n18539), .B2(n19372), .ZN(
        n1732) );
  OAI221_X1 U2256 ( .B1(n19619), .B2(n18550), .C1(n19651), .C2(n18547), .A(
        n1714), .ZN(n1711) );
  AOI22_X1 U2257 ( .A1(n18544), .A2(n17754), .B1(n18539), .B2(n19371), .ZN(
        n1714) );
  OAI221_X1 U2258 ( .B1(n19618), .B2(n18550), .C1(n19650), .C2(n18547), .A(
        n1696), .ZN(n1693) );
  AOI22_X1 U2259 ( .A1(n18544), .A2(n17755), .B1(n18539), .B2(n19370), .ZN(
        n1696) );
  OAI221_X1 U2260 ( .B1(n19617), .B2(n18550), .C1(n19649), .C2(n18547), .A(
        n1678), .ZN(n1675) );
  AOI22_X1 U2261 ( .A1(n18544), .A2(n17756), .B1(n18539), .B2(n19369), .ZN(
        n1678) );
  OAI221_X1 U2262 ( .B1(n19616), .B2(n18550), .C1(n19648), .C2(n18547), .A(
        n1660), .ZN(n1657) );
  AOI22_X1 U2263 ( .A1(n18544), .A2(n17757), .B1(n18539), .B2(n19368), .ZN(
        n1660) );
  OAI221_X1 U2264 ( .B1(n19615), .B2(n18550), .C1(n19647), .C2(n18547), .A(
        n1632), .ZN(n1623) );
  AOI22_X1 U2265 ( .A1(n18544), .A2(n17758), .B1(n18539), .B2(n19367), .ZN(
        n1632) );
  OAI22_X1 U2266 ( .A1(n18513), .A2(n18806), .B1(n17871), .B2(n18815), .ZN(
        n3198) );
  OAI22_X1 U2267 ( .A1(n18510), .A2(n18806), .B1(n17872), .B2(n18815), .ZN(
        n3199) );
  OAI22_X1 U2268 ( .A1(n18507), .A2(n18806), .B1(n17873), .B2(n18815), .ZN(
        n3200) );
  OAI22_X1 U2269 ( .A1(n18504), .A2(n18806), .B1(n17874), .B2(n18815), .ZN(
        n3201) );
  OAI22_X1 U2270 ( .A1(n18501), .A2(n18806), .B1(n17875), .B2(n18814), .ZN(
        n3202) );
  OAI22_X1 U2271 ( .A1(n18498), .A2(n18806), .B1(n17876), .B2(n18814), .ZN(
        n3203) );
  OAI22_X1 U2272 ( .A1(n18492), .A2(n18806), .B1(n17878), .B2(n18814), .ZN(
        n3205) );
  OAI22_X1 U2273 ( .A1(n18489), .A2(n18806), .B1(n17879), .B2(n18813), .ZN(
        n3206) );
  OAI22_X1 U2274 ( .A1(n18486), .A2(n18806), .B1(n17880), .B2(n18813), .ZN(
        n3207) );
  OAI22_X1 U2275 ( .A1(n18483), .A2(n18806), .B1(n17881), .B2(n18813), .ZN(
        n3208) );
  OAI22_X1 U2276 ( .A1(n18480), .A2(n18806), .B1(n17882), .B2(n18813), .ZN(
        n3209) );
  OAI22_X1 U2277 ( .A1(n18477), .A2(n18807), .B1(n17883), .B2(n18812), .ZN(
        n3210) );
  OAI22_X1 U2278 ( .A1(n18474), .A2(n18807), .B1(n17884), .B2(n18812), .ZN(
        n3211) );
  OAI22_X1 U2279 ( .A1(n18471), .A2(n18807), .B1(n17885), .B2(n18812), .ZN(
        n3212) );
  OAI22_X1 U2280 ( .A1(n18468), .A2(n18807), .B1(n17886), .B2(n18812), .ZN(
        n3213) );
  OAI22_X1 U2281 ( .A1(n18465), .A2(n18807), .B1(n17887), .B2(n18811), .ZN(
        n3214) );
  OAI22_X1 U2282 ( .A1(n18462), .A2(n18807), .B1(n17888), .B2(n18811), .ZN(
        n3215) );
  OAI22_X1 U2283 ( .A1(n18459), .A2(n18807), .B1(n17889), .B2(n18811), .ZN(
        n3216) );
  OAI22_X1 U2284 ( .A1(n18456), .A2(n18807), .B1(n17890), .B2(n18811), .ZN(
        n3217) );
  OAI22_X1 U2285 ( .A1(n18453), .A2(n18807), .B1(n17891), .B2(n18810), .ZN(
        n3218) );
  OAI22_X1 U2286 ( .A1(n18450), .A2(n18807), .B1(n17892), .B2(n18810), .ZN(
        n3219) );
  OAI22_X1 U2287 ( .A1(n18447), .A2(n18807), .B1(n17893), .B2(n18810), .ZN(
        n3220) );
  OAI22_X1 U2288 ( .A1(n18444), .A2(n18807), .B1(n17894), .B2(n18810), .ZN(
        n3221) );
  OAI22_X1 U2289 ( .A1(n18488), .A2(n18972), .B1(n18075), .B2(n18975), .ZN(
        n3829) );
  OAI22_X1 U2290 ( .A1(n18485), .A2(n18972), .B1(n18076), .B2(n18975), .ZN(
        n3813) );
  OAI22_X1 U2291 ( .A1(n18482), .A2(n18972), .B1(n18077), .B2(n18975), .ZN(
        n3797) );
  OAI22_X1 U2292 ( .A1(n18479), .A2(n18972), .B1(n18078), .B2(n18975), .ZN(
        n3781) );
  OAI22_X1 U2293 ( .A1(n18476), .A2(n18972), .B1(n18079), .B2(n18976), .ZN(
        n3765) );
  OAI22_X1 U2294 ( .A1(n18473), .A2(n18972), .B1(n18080), .B2(n18976), .ZN(
        n3749) );
  OAI22_X1 U2295 ( .A1(n18470), .A2(n18972), .B1(n18081), .B2(n18976), .ZN(
        n3733) );
  OAI22_X1 U2296 ( .A1(n18467), .A2(n18972), .B1(n18082), .B2(n18976), .ZN(
        n3717) );
  OAI22_X1 U2297 ( .A1(n18464), .A2(n18972), .B1(n18083), .B2(n18977), .ZN(
        n3701) );
  OAI22_X1 U2298 ( .A1(n18461), .A2(n18972), .B1(n18084), .B2(n18977), .ZN(
        n3685) );
  OAI22_X1 U2299 ( .A1(n18458), .A2(n18972), .B1(n18085), .B2(n18977), .ZN(
        n3669) );
  OAI22_X1 U2300 ( .A1(n18455), .A2(n18972), .B1(n18086), .B2(n18977), .ZN(
        n3653) );
  OAI22_X1 U2301 ( .A1(n18452), .A2(n18971), .B1(n18087), .B2(n18978), .ZN(
        n3637) );
  OAI22_X1 U2302 ( .A1(n18449), .A2(n18971), .B1(n18088), .B2(n18978), .ZN(
        n3621) );
  OAI22_X1 U2303 ( .A1(n18446), .A2(n18971), .B1(n18089), .B2(n18978), .ZN(
        n3605) );
  OAI22_X1 U2304 ( .A1(n18443), .A2(n18971), .B1(n18090), .B2(n18978), .ZN(
        n3589) );
  OAI22_X1 U2305 ( .A1(n18440), .A2(n18971), .B1(n18091), .B2(n18979), .ZN(
        n3573) );
  OAI22_X1 U2306 ( .A1(n18437), .A2(n18971), .B1(n18092), .B2(n18979), .ZN(
        n3557) );
  OAI22_X1 U2307 ( .A1(n18434), .A2(n18971), .B1(n18093), .B2(n18979), .ZN(
        n3541) );
  OAI22_X1 U2308 ( .A1(n18431), .A2(n18971), .B1(n18094), .B2(n18979), .ZN(
        n3525) );
  OAI22_X1 U2309 ( .A1(n18428), .A2(n18971), .B1(n18095), .B2(n18980), .ZN(
        n3509) );
  OAI22_X1 U2310 ( .A1(n18425), .A2(n18971), .B1(n18096), .B2(n18980), .ZN(
        n3493) );
  OAI22_X1 U2311 ( .A1(n18422), .A2(n18971), .B1(n18097), .B2(n18980), .ZN(
        n3477) );
  OAI22_X1 U2312 ( .A1(n18419), .A2(n18971), .B1(n18098), .B2(n18980), .ZN(
        n3461) );
  OAI22_X1 U2313 ( .A1(n18513), .A2(n18872), .B1(n18099), .B2(n18881), .ZN(
        n3390) );
  OAI22_X1 U2314 ( .A1(n18510), .A2(n18872), .B1(n18100), .B2(n18881), .ZN(
        n3391) );
  OAI22_X1 U2315 ( .A1(n18507), .A2(n18872), .B1(n18101), .B2(n18881), .ZN(
        n3392) );
  OAI22_X1 U2316 ( .A1(n18504), .A2(n18872), .B1(n18102), .B2(n18881), .ZN(
        n3393) );
  OAI22_X1 U2317 ( .A1(n18501), .A2(n18872), .B1(n18103), .B2(n18880), .ZN(
        n3394) );
  OAI22_X1 U2318 ( .A1(n18498), .A2(n18872), .B1(n18104), .B2(n18880), .ZN(
        n3395) );
  OAI22_X1 U2319 ( .A1(n18495), .A2(n18872), .B1(n18105), .B2(n18880), .ZN(
        n3396) );
  OAI22_X1 U2320 ( .A1(n18492), .A2(n18872), .B1(n18106), .B2(n18880), .ZN(
        n3397) );
  OAI22_X1 U2321 ( .A1(n18489), .A2(n18872), .B1(n18107), .B2(n18879), .ZN(
        n3398) );
  OAI22_X1 U2322 ( .A1(n18486), .A2(n18872), .B1(n18108), .B2(n18879), .ZN(
        n3399) );
  OAI22_X1 U2323 ( .A1(n18483), .A2(n18872), .B1(n18109), .B2(n18879), .ZN(
        n3400) );
  OAI22_X1 U2324 ( .A1(n18480), .A2(n18872), .B1(n18110), .B2(n18879), .ZN(
        n3401) );
  OAI22_X1 U2325 ( .A1(n18477), .A2(n18873), .B1(n18111), .B2(n18878), .ZN(
        n3402) );
  OAI22_X1 U2326 ( .A1(n18474), .A2(n18873), .B1(n18112), .B2(n18878), .ZN(
        n3403) );
  OAI22_X1 U2327 ( .A1(n18471), .A2(n18873), .B1(n18113), .B2(n18878), .ZN(
        n3404) );
  OAI22_X1 U2328 ( .A1(n18468), .A2(n18873), .B1(n18114), .B2(n18878), .ZN(
        n3405) );
  OAI22_X1 U2329 ( .A1(n18465), .A2(n18873), .B1(n18115), .B2(n18877), .ZN(
        n3406) );
  OAI22_X1 U2330 ( .A1(n18462), .A2(n18873), .B1(n18116), .B2(n18877), .ZN(
        n3407) );
  OAI22_X1 U2331 ( .A1(n18459), .A2(n18873), .B1(n18117), .B2(n18877), .ZN(
        n3408) );
  OAI22_X1 U2332 ( .A1(n18456), .A2(n18873), .B1(n18118), .B2(n18877), .ZN(
        n3409) );
  OAI22_X1 U2333 ( .A1(n18453), .A2(n18873), .B1(n18119), .B2(n18876), .ZN(
        n3410) );
  OAI22_X1 U2334 ( .A1(n18450), .A2(n18873), .B1(n18120), .B2(n18876), .ZN(
        n3411) );
  OAI22_X1 U2335 ( .A1(n18447), .A2(n18873), .B1(n18121), .B2(n18876), .ZN(
        n3412) );
  OAI22_X1 U2336 ( .A1(n18444), .A2(n18873), .B1(n18122), .B2(n18876), .ZN(
        n3413) );
  OAI22_X1 U2337 ( .A1(n18441), .A2(n18806), .B1(n18219), .B2(n18809), .ZN(
        n3222) );
  OAI22_X1 U2338 ( .A1(n18438), .A2(n18807), .B1(n18220), .B2(n18809), .ZN(
        n3223) );
  OAI22_X1 U2339 ( .A1(n18435), .A2(n18806), .B1(n18221), .B2(n18809), .ZN(
        n3224) );
  OAI22_X1 U2340 ( .A1(n18432), .A2(n18807), .B1(n18222), .B2(n18809), .ZN(
        n3225) );
  OAI22_X1 U2341 ( .A1(n18429), .A2(n18806), .B1(n18223), .B2(n18808), .ZN(
        n3226) );
  OAI22_X1 U2342 ( .A1(n18426), .A2(n18807), .B1(n18224), .B2(n18808), .ZN(
        n3227) );
  OAI22_X1 U2343 ( .A1(n18423), .A2(n18806), .B1(n18225), .B2(n18808), .ZN(
        n3228) );
  OAI22_X1 U2344 ( .A1(n18420), .A2(n18807), .B1(n18226), .B2(n18808), .ZN(
        n3229) );
  OAI22_X1 U2345 ( .A1(n18512), .A2(n18972), .B1(n18283), .B2(n18973), .ZN(
        n3957) );
  OAI22_X1 U2346 ( .A1(n18509), .A2(n18971), .B1(n18284), .B2(n18973), .ZN(
        n3941) );
  OAI22_X1 U2347 ( .A1(n18506), .A2(n18972), .B1(n18285), .B2(n18973), .ZN(
        n3925) );
  OAI22_X1 U2348 ( .A1(n18503), .A2(n18971), .B1(n18286), .B2(n18973), .ZN(
        n3909) );
  OAI22_X1 U2349 ( .A1(n18500), .A2(n18972), .B1(n18287), .B2(n18974), .ZN(
        n3893) );
  OAI22_X1 U2350 ( .A1(n18497), .A2(n18971), .B1(n18288), .B2(n18974), .ZN(
        n3877) );
  OAI22_X1 U2351 ( .A1(n18494), .A2(n18972), .B1(n18289), .B2(n18974), .ZN(
        n3861) );
  OAI22_X1 U2352 ( .A1(n18491), .A2(n18971), .B1(n18290), .B2(n18974), .ZN(
        n3845) );
  OAI22_X1 U2353 ( .A1(n18441), .A2(n18872), .B1(n18291), .B2(n18875), .ZN(
        n3414) );
  OAI22_X1 U2354 ( .A1(n18438), .A2(n18873), .B1(n18292), .B2(n18875), .ZN(
        n3415) );
  OAI22_X1 U2355 ( .A1(n18435), .A2(n18872), .B1(n18293), .B2(n18875), .ZN(
        n3416) );
  OAI22_X1 U2356 ( .A1(n18432), .A2(n18873), .B1(n18294), .B2(n18875), .ZN(
        n3417) );
  OAI22_X1 U2357 ( .A1(n18429), .A2(n18872), .B1(n18295), .B2(n18874), .ZN(
        n3418) );
  OAI22_X1 U2358 ( .A1(n18426), .A2(n18873), .B1(n18296), .B2(n18874), .ZN(
        n3419) );
  OAI22_X1 U2359 ( .A1(n18423), .A2(n18872), .B1(n18297), .B2(n18874), .ZN(
        n3420) );
  OAI22_X1 U2360 ( .A1(n18420), .A2(n18873), .B1(n18298), .B2(n18874), .ZN(
        n3421) );
  OAI22_X1 U2361 ( .A1(n18513), .A2(n18784), .B1(n17791), .B2(n18793), .ZN(
        n3134) );
  OAI22_X1 U2362 ( .A1(n18510), .A2(n18784), .B1(n17792), .B2(n18793), .ZN(
        n3135) );
  OAI22_X1 U2363 ( .A1(n18507), .A2(n18784), .B1(n17793), .B2(n18793), .ZN(
        n3136) );
  OAI22_X1 U2364 ( .A1(n18504), .A2(n18784), .B1(n17794), .B2(n18793), .ZN(
        n3137) );
  OAI22_X1 U2365 ( .A1(n18501), .A2(n18784), .B1(n17795), .B2(n18792), .ZN(
        n3138) );
  OAI22_X1 U2366 ( .A1(n18498), .A2(n18784), .B1(n17796), .B2(n18792), .ZN(
        n3139) );
  OAI22_X1 U2367 ( .A1(n18495), .A2(n18784), .B1(n17797), .B2(n18792), .ZN(
        n3140) );
  OAI22_X1 U2368 ( .A1(n18492), .A2(n18784), .B1(n17798), .B2(n18792), .ZN(
        n3141) );
  OAI22_X1 U2369 ( .A1(n18489), .A2(n18784), .B1(n17799), .B2(n18791), .ZN(
        n3142) );
  OAI22_X1 U2370 ( .A1(n18486), .A2(n18784), .B1(n17800), .B2(n18791), .ZN(
        n3143) );
  OAI22_X1 U2371 ( .A1(n18483), .A2(n18784), .B1(n17801), .B2(n18791), .ZN(
        n3144) );
  OAI22_X1 U2372 ( .A1(n18480), .A2(n18784), .B1(n17802), .B2(n18791), .ZN(
        n3145) );
  OAI22_X1 U2373 ( .A1(n18477), .A2(n18785), .B1(n17803), .B2(n18790), .ZN(
        n3146) );
  OAI22_X1 U2374 ( .A1(n18474), .A2(n18785), .B1(n17804), .B2(n18790), .ZN(
        n3147) );
  OAI22_X1 U2375 ( .A1(n18471), .A2(n18785), .B1(n17805), .B2(n18790), .ZN(
        n3148) );
  OAI22_X1 U2376 ( .A1(n18468), .A2(n18785), .B1(n17806), .B2(n18790), .ZN(
        n3149) );
  OAI22_X1 U2377 ( .A1(n18465), .A2(n18785), .B1(n17807), .B2(n18789), .ZN(
        n3150) );
  OAI22_X1 U2378 ( .A1(n18462), .A2(n18785), .B1(n17808), .B2(n18789), .ZN(
        n3151) );
  OAI22_X1 U2379 ( .A1(n18459), .A2(n18785), .B1(n17809), .B2(n18789), .ZN(
        n3152) );
  OAI22_X1 U2380 ( .A1(n18456), .A2(n18785), .B1(n17810), .B2(n18789), .ZN(
        n3153) );
  OAI22_X1 U2381 ( .A1(n18453), .A2(n18785), .B1(n17811), .B2(n18788), .ZN(
        n3154) );
  OAI22_X1 U2382 ( .A1(n18450), .A2(n18785), .B1(n17812), .B2(n18788), .ZN(
        n3155) );
  OAI22_X1 U2383 ( .A1(n18447), .A2(n18785), .B1(n17813), .B2(n18788), .ZN(
        n3156) );
  OAI22_X1 U2384 ( .A1(n18444), .A2(n18785), .B1(n17814), .B2(n18788), .ZN(
        n3157) );
  OAI22_X1 U2385 ( .A1(n18513), .A2(n18850), .B1(n17847), .B2(n18859), .ZN(
        n3326) );
  OAI22_X1 U2386 ( .A1(n18510), .A2(n18850), .B1(n17848), .B2(n18859), .ZN(
        n3327) );
  OAI22_X1 U2387 ( .A1(n18507), .A2(n18850), .B1(n17849), .B2(n18859), .ZN(
        n3328) );
  OAI22_X1 U2388 ( .A1(n18504), .A2(n18850), .B1(n17850), .B2(n18859), .ZN(
        n3329) );
  OAI22_X1 U2389 ( .A1(n18501), .A2(n18850), .B1(n17851), .B2(n18858), .ZN(
        n3330) );
  OAI22_X1 U2390 ( .A1(n18498), .A2(n18850), .B1(n17852), .B2(n18858), .ZN(
        n3331) );
  OAI22_X1 U2391 ( .A1(n18495), .A2(n18850), .B1(n17853), .B2(n18858), .ZN(
        n3332) );
  OAI22_X1 U2392 ( .A1(n18492), .A2(n18850), .B1(n17854), .B2(n18858), .ZN(
        n3333) );
  OAI22_X1 U2393 ( .A1(n18489), .A2(n18850), .B1(n17855), .B2(n18857), .ZN(
        n3334) );
  OAI22_X1 U2394 ( .A1(n18486), .A2(n18850), .B1(n17856), .B2(n18857), .ZN(
        n3335) );
  OAI22_X1 U2395 ( .A1(n18483), .A2(n18850), .B1(n17857), .B2(n18857), .ZN(
        n3336) );
  OAI22_X1 U2396 ( .A1(n18480), .A2(n18850), .B1(n17858), .B2(n18857), .ZN(
        n3337) );
  OAI22_X1 U2397 ( .A1(n18477), .A2(n18851), .B1(n17859), .B2(n18856), .ZN(
        n3338) );
  OAI22_X1 U2398 ( .A1(n18474), .A2(n18851), .B1(n17860), .B2(n18856), .ZN(
        n3339) );
  OAI22_X1 U2399 ( .A1(n18471), .A2(n18851), .B1(n17861), .B2(n18856), .ZN(
        n3340) );
  OAI22_X1 U2400 ( .A1(n18468), .A2(n18851), .B1(n17862), .B2(n18856), .ZN(
        n3341) );
  OAI22_X1 U2401 ( .A1(n18465), .A2(n18851), .B1(n17863), .B2(n18855), .ZN(
        n3342) );
  OAI22_X1 U2402 ( .A1(n18462), .A2(n18851), .B1(n17864), .B2(n18855), .ZN(
        n3343) );
  OAI22_X1 U2403 ( .A1(n18459), .A2(n18851), .B1(n17865), .B2(n18855), .ZN(
        n3344) );
  OAI22_X1 U2404 ( .A1(n18456), .A2(n18851), .B1(n17866), .B2(n18855), .ZN(
        n3345) );
  OAI22_X1 U2405 ( .A1(n18453), .A2(n18851), .B1(n17867), .B2(n18854), .ZN(
        n3346) );
  OAI22_X1 U2406 ( .A1(n18450), .A2(n18851), .B1(n17868), .B2(n18854), .ZN(
        n3347) );
  OAI22_X1 U2407 ( .A1(n18447), .A2(n18851), .B1(n17869), .B2(n18854), .ZN(
        n3348) );
  OAI22_X1 U2408 ( .A1(n18444), .A2(n18851), .B1(n17870), .B2(n18854), .ZN(
        n3349) );
  OAI22_X1 U2409 ( .A1(n18441), .A2(n18784), .B1(n18195), .B2(n18787), .ZN(
        n3158) );
  OAI22_X1 U2410 ( .A1(n18438), .A2(n18785), .B1(n18196), .B2(n18787), .ZN(
        n3159) );
  OAI22_X1 U2411 ( .A1(n18435), .A2(n18784), .B1(n18197), .B2(n18787), .ZN(
        n3160) );
  OAI22_X1 U2412 ( .A1(n18432), .A2(n18785), .B1(n18198), .B2(n18787), .ZN(
        n3161) );
  OAI22_X1 U2413 ( .A1(n18429), .A2(n18784), .B1(n18199), .B2(n18786), .ZN(
        n3162) );
  OAI22_X1 U2414 ( .A1(n18426), .A2(n18785), .B1(n18200), .B2(n18786), .ZN(
        n3163) );
  OAI22_X1 U2415 ( .A1(n18423), .A2(n18784), .B1(n18201), .B2(n18786), .ZN(
        n3164) );
  OAI22_X1 U2416 ( .A1(n18420), .A2(n18785), .B1(n18202), .B2(n18786), .ZN(
        n3165) );
  OAI22_X1 U2417 ( .A1(n18441), .A2(n18850), .B1(n18211), .B2(n18853), .ZN(
        n3350) );
  OAI22_X1 U2418 ( .A1(n18438), .A2(n18851), .B1(n18212), .B2(n18853), .ZN(
        n3351) );
  OAI22_X1 U2419 ( .A1(n18435), .A2(n18850), .B1(n18213), .B2(n18853), .ZN(
        n3352) );
  OAI22_X1 U2420 ( .A1(n18432), .A2(n18851), .B1(n18214), .B2(n18853), .ZN(
        n3353) );
  OAI22_X1 U2421 ( .A1(n18429), .A2(n18850), .B1(n18215), .B2(n18852), .ZN(
        n3354) );
  OAI22_X1 U2422 ( .A1(n18426), .A2(n18851), .B1(n18216), .B2(n18852), .ZN(
        n3355) );
  OAI22_X1 U2423 ( .A1(n18423), .A2(n18850), .B1(n18217), .B2(n18852), .ZN(
        n3356) );
  OAI22_X1 U2424 ( .A1(n18420), .A2(n18851), .B1(n18218), .B2(n18852), .ZN(
        n3357) );
  OAI22_X1 U2425 ( .A1(n19054), .A2(n18512), .B1(n2496), .B2(n19046), .ZN(
        n9174) );
  OAI22_X1 U2426 ( .A1(n19054), .A2(n18509), .B1(n2487), .B2(n19046), .ZN(
        n9175) );
  OAI22_X1 U2427 ( .A1(n19053), .A2(n18506), .B1(n2478), .B2(n19046), .ZN(
        n9176) );
  OAI22_X1 U2428 ( .A1(n19053), .A2(n18503), .B1(n2469), .B2(n19046), .ZN(
        n9177) );
  OAI22_X1 U2429 ( .A1(n19053), .A2(n18500), .B1(n2460), .B2(n19046), .ZN(
        n9178) );
  OAI22_X1 U2430 ( .A1(n19053), .A2(n18497), .B1(n2451), .B2(n19046), .ZN(
        n9179) );
  OAI22_X1 U2431 ( .A1(n19053), .A2(n18494), .B1(n2442), .B2(n19046), .ZN(
        n9180) );
  OAI22_X1 U2432 ( .A1(n19052), .A2(n18491), .B1(n2433), .B2(n19046), .ZN(
        n9181) );
  OAI22_X1 U2433 ( .A1(n19052), .A2(n18488), .B1(n2424), .B2(n19046), .ZN(
        n9182) );
  OAI22_X1 U2434 ( .A1(n19052), .A2(n18485), .B1(n2415), .B2(n19046), .ZN(
        n9183) );
  OAI22_X1 U2435 ( .A1(n19052), .A2(n18482), .B1(n2406), .B2(n19046), .ZN(
        n9184) );
  OAI22_X1 U2436 ( .A1(n19052), .A2(n18479), .B1(n2397), .B2(n19046), .ZN(
        n9185) );
  OAI22_X1 U2437 ( .A1(n19051), .A2(n18476), .B1(n2388), .B2(n19047), .ZN(
        n9186) );
  OAI22_X1 U2438 ( .A1(n19051), .A2(n18473), .B1(n2379), .B2(n19047), .ZN(
        n9187) );
  OAI22_X1 U2439 ( .A1(n19051), .A2(n18470), .B1(n2370), .B2(n19047), .ZN(
        n9188) );
  OAI22_X1 U2440 ( .A1(n19051), .A2(n18467), .B1(n2361), .B2(n19047), .ZN(
        n9189) );
  OAI22_X1 U2441 ( .A1(n19051), .A2(n18464), .B1(n2352), .B2(n19047), .ZN(
        n9190) );
  OAI22_X1 U2442 ( .A1(n19050), .A2(n18461), .B1(n2343), .B2(n19047), .ZN(
        n9191) );
  OAI22_X1 U2443 ( .A1(n19050), .A2(n18458), .B1(n2334), .B2(n19047), .ZN(
        n9192) );
  OAI22_X1 U2444 ( .A1(n19050), .A2(n18455), .B1(n2325), .B2(n19047), .ZN(
        n9193) );
  OAI22_X1 U2445 ( .A1(n19050), .A2(n18452), .B1(n2316), .B2(n19047), .ZN(
        n9194) );
  OAI22_X1 U2446 ( .A1(n19050), .A2(n18449), .B1(n2307), .B2(n19047), .ZN(
        n9195) );
  OAI22_X1 U2447 ( .A1(n19049), .A2(n18446), .B1(n2298), .B2(n19047), .ZN(
        n9196) );
  OAI22_X1 U2448 ( .A1(n19049), .A2(n18443), .B1(n2289), .B2(n19047), .ZN(
        n9197) );
  OAI22_X1 U2449 ( .A1(n18513), .A2(n18762), .B1(n17895), .B2(n18771), .ZN(
        n3070) );
  OAI22_X1 U2450 ( .A1(n18510), .A2(n18762), .B1(n17896), .B2(n18771), .ZN(
        n3071) );
  OAI22_X1 U2451 ( .A1(n18507), .A2(n18762), .B1(n17897), .B2(n18771), .ZN(
        n3072) );
  OAI22_X1 U2452 ( .A1(n18504), .A2(n18762), .B1(n17898), .B2(n18771), .ZN(
        n3073) );
  OAI22_X1 U2453 ( .A1(n18501), .A2(n18762), .B1(n17899), .B2(n18770), .ZN(
        n3074) );
  OAI22_X1 U2454 ( .A1(n18498), .A2(n18762), .B1(n17900), .B2(n18770), .ZN(
        n3075) );
  OAI22_X1 U2455 ( .A1(n18495), .A2(n18762), .B1(n17901), .B2(n18770), .ZN(
        n3076) );
  OAI22_X1 U2456 ( .A1(n18492), .A2(n18762), .B1(n17902), .B2(n18770), .ZN(
        n3077) );
  OAI22_X1 U2457 ( .A1(n18489), .A2(n18762), .B1(n17903), .B2(n18769), .ZN(
        n3078) );
  OAI22_X1 U2458 ( .A1(n18486), .A2(n18762), .B1(n17904), .B2(n18769), .ZN(
        n3079) );
  OAI22_X1 U2459 ( .A1(n18483), .A2(n18762), .B1(n17905), .B2(n18769), .ZN(
        n3080) );
  OAI22_X1 U2460 ( .A1(n18480), .A2(n18762), .B1(n17906), .B2(n18769), .ZN(
        n3081) );
  OAI22_X1 U2461 ( .A1(n18477), .A2(n18763), .B1(n17907), .B2(n18768), .ZN(
        n3082) );
  OAI22_X1 U2462 ( .A1(n18474), .A2(n18763), .B1(n17908), .B2(n18768), .ZN(
        n3083) );
  OAI22_X1 U2463 ( .A1(n18471), .A2(n18763), .B1(n17909), .B2(n18768), .ZN(
        n3084) );
  OAI22_X1 U2464 ( .A1(n18468), .A2(n18763), .B1(n17910), .B2(n18768), .ZN(
        n3085) );
  OAI22_X1 U2465 ( .A1(n18465), .A2(n18763), .B1(n17911), .B2(n18767), .ZN(
        n3086) );
  OAI22_X1 U2466 ( .A1(n18462), .A2(n18763), .B1(n17912), .B2(n18767), .ZN(
        n3087) );
  OAI22_X1 U2467 ( .A1(n18459), .A2(n18763), .B1(n17913), .B2(n18767), .ZN(
        n3088) );
  OAI22_X1 U2468 ( .A1(n18456), .A2(n18763), .B1(n17914), .B2(n18767), .ZN(
        n3089) );
  OAI22_X1 U2469 ( .A1(n18453), .A2(n18763), .B1(n17915), .B2(n18766), .ZN(
        n3090) );
  OAI22_X1 U2470 ( .A1(n18450), .A2(n18763), .B1(n17916), .B2(n18766), .ZN(
        n3091) );
  OAI22_X1 U2471 ( .A1(n18447), .A2(n18763), .B1(n17917), .B2(n18766), .ZN(
        n3092) );
  OAI22_X1 U2472 ( .A1(n18444), .A2(n18763), .B1(n17918), .B2(n18766), .ZN(
        n3093) );
  OAI22_X1 U2473 ( .A1(n18513), .A2(n18839), .B1(n18123), .B2(n18848), .ZN(
        n3294) );
  OAI22_X1 U2474 ( .A1(n18510), .A2(n18839), .B1(n18124), .B2(n18848), .ZN(
        n3295) );
  OAI22_X1 U2475 ( .A1(n18507), .A2(n18839), .B1(n18125), .B2(n18848), .ZN(
        n3296) );
  OAI22_X1 U2476 ( .A1(n18504), .A2(n18839), .B1(n18126), .B2(n18848), .ZN(
        n3297) );
  OAI22_X1 U2477 ( .A1(n18501), .A2(n18839), .B1(n18127), .B2(n18847), .ZN(
        n3298) );
  OAI22_X1 U2478 ( .A1(n18498), .A2(n18839), .B1(n18128), .B2(n18847), .ZN(
        n3299) );
  OAI22_X1 U2479 ( .A1(n18495), .A2(n18839), .B1(n18129), .B2(n18847), .ZN(
        n3300) );
  OAI22_X1 U2480 ( .A1(n18492), .A2(n18839), .B1(n18130), .B2(n18847), .ZN(
        n3301) );
  OAI22_X1 U2481 ( .A1(n18489), .A2(n18839), .B1(n18131), .B2(n18846), .ZN(
        n3302) );
  OAI22_X1 U2482 ( .A1(n18486), .A2(n18839), .B1(n18132), .B2(n18846), .ZN(
        n3303) );
  OAI22_X1 U2483 ( .A1(n18483), .A2(n18839), .B1(n18133), .B2(n18846), .ZN(
        n3304) );
  OAI22_X1 U2484 ( .A1(n18480), .A2(n18839), .B1(n18134), .B2(n18846), .ZN(
        n3305) );
  OAI22_X1 U2485 ( .A1(n18477), .A2(n18840), .B1(n18135), .B2(n18845), .ZN(
        n3306) );
  OAI22_X1 U2486 ( .A1(n18474), .A2(n18840), .B1(n18136), .B2(n18845), .ZN(
        n3307) );
  OAI22_X1 U2487 ( .A1(n18471), .A2(n18840), .B1(n18137), .B2(n18845), .ZN(
        n3308) );
  OAI22_X1 U2488 ( .A1(n18468), .A2(n18840), .B1(n18138), .B2(n18845), .ZN(
        n3309) );
  OAI22_X1 U2489 ( .A1(n18465), .A2(n18840), .B1(n18139), .B2(n18844), .ZN(
        n3310) );
  OAI22_X1 U2490 ( .A1(n18462), .A2(n18840), .B1(n18140), .B2(n18844), .ZN(
        n3311) );
  OAI22_X1 U2491 ( .A1(n18459), .A2(n18840), .B1(n18141), .B2(n18844), .ZN(
        n3312) );
  OAI22_X1 U2492 ( .A1(n18456), .A2(n18840), .B1(n18142), .B2(n18844), .ZN(
        n3313) );
  OAI22_X1 U2493 ( .A1(n18453), .A2(n18840), .B1(n18143), .B2(n18843), .ZN(
        n3314) );
  OAI22_X1 U2494 ( .A1(n18450), .A2(n18840), .B1(n18144), .B2(n18843), .ZN(
        n3315) );
  OAI22_X1 U2495 ( .A1(n18447), .A2(n18840), .B1(n18145), .B2(n18843), .ZN(
        n3316) );
  OAI22_X1 U2496 ( .A1(n18444), .A2(n18840), .B1(n18146), .B2(n18843), .ZN(
        n3317) );
  OAI22_X1 U2497 ( .A1(n18441), .A2(n18762), .B1(n18227), .B2(n18765), .ZN(
        n3094) );
  OAI22_X1 U2498 ( .A1(n18438), .A2(n18763), .B1(n18228), .B2(n18765), .ZN(
        n3095) );
  OAI22_X1 U2499 ( .A1(n18435), .A2(n18762), .B1(n18229), .B2(n18765), .ZN(
        n3096) );
  OAI22_X1 U2500 ( .A1(n18432), .A2(n18763), .B1(n18230), .B2(n18765), .ZN(
        n3097) );
  OAI22_X1 U2501 ( .A1(n18429), .A2(n18762), .B1(n18231), .B2(n18764), .ZN(
        n3098) );
  OAI22_X1 U2502 ( .A1(n18426), .A2(n18763), .B1(n18232), .B2(n18764), .ZN(
        n3099) );
  OAI22_X1 U2503 ( .A1(n18423), .A2(n18762), .B1(n18233), .B2(n18764), .ZN(
        n3100) );
  OAI22_X1 U2504 ( .A1(n18420), .A2(n18763), .B1(n18234), .B2(n18764), .ZN(
        n3101) );
  OAI22_X1 U2505 ( .A1(n18441), .A2(n18839), .B1(n18299), .B2(n18842), .ZN(
        n3318) );
  OAI22_X1 U2506 ( .A1(n18438), .A2(n18840), .B1(n18300), .B2(n18842), .ZN(
        n3319) );
  OAI22_X1 U2507 ( .A1(n18435), .A2(n18839), .B1(n18301), .B2(n18842), .ZN(
        n3320) );
  OAI22_X1 U2508 ( .A1(n18432), .A2(n18840), .B1(n18302), .B2(n18842), .ZN(
        n3321) );
  OAI22_X1 U2509 ( .A1(n18429), .A2(n18839), .B1(n18303), .B2(n18841), .ZN(
        n3322) );
  OAI22_X1 U2510 ( .A1(n18426), .A2(n18840), .B1(n18304), .B2(n18841), .ZN(
        n3323) );
  OAI22_X1 U2511 ( .A1(n18423), .A2(n18839), .B1(n18305), .B2(n18841), .ZN(
        n3324) );
  OAI22_X1 U2512 ( .A1(n18420), .A2(n18840), .B1(n18306), .B2(n18841), .ZN(
        n3325) );
  OAI22_X1 U2513 ( .A1(n18514), .A2(n18751), .B1(n17815), .B2(n18760), .ZN(
        n3038) );
  OAI22_X1 U2514 ( .A1(n18511), .A2(n18751), .B1(n17816), .B2(n18760), .ZN(
        n3039) );
  OAI22_X1 U2515 ( .A1(n18508), .A2(n18751), .B1(n17817), .B2(n18760), .ZN(
        n3040) );
  OAI22_X1 U2516 ( .A1(n18505), .A2(n18751), .B1(n17818), .B2(n18760), .ZN(
        n3041) );
  OAI22_X1 U2517 ( .A1(n18502), .A2(n18751), .B1(n17819), .B2(n18759), .ZN(
        n3042) );
  OAI22_X1 U2518 ( .A1(n18499), .A2(n18751), .B1(n17820), .B2(n18759), .ZN(
        n3043) );
  OAI22_X1 U2519 ( .A1(n18496), .A2(n18751), .B1(n17821), .B2(n18759), .ZN(
        n3044) );
  OAI22_X1 U2520 ( .A1(n18493), .A2(n18751), .B1(n17822), .B2(n18759), .ZN(
        n3045) );
  OAI22_X1 U2521 ( .A1(n18490), .A2(n18751), .B1(n17823), .B2(n18758), .ZN(
        n3046) );
  OAI22_X1 U2522 ( .A1(n18487), .A2(n18751), .B1(n17824), .B2(n18758), .ZN(
        n3047) );
  OAI22_X1 U2523 ( .A1(n18484), .A2(n18751), .B1(n17825), .B2(n18758), .ZN(
        n3048) );
  OAI22_X1 U2524 ( .A1(n18481), .A2(n18751), .B1(n17826), .B2(n18758), .ZN(
        n3049) );
  OAI22_X1 U2525 ( .A1(n18478), .A2(n18752), .B1(n17827), .B2(n18757), .ZN(
        n3050) );
  OAI22_X1 U2526 ( .A1(n18475), .A2(n18752), .B1(n17828), .B2(n18757), .ZN(
        n3051) );
  OAI22_X1 U2527 ( .A1(n18472), .A2(n18752), .B1(n17829), .B2(n18757), .ZN(
        n3052) );
  OAI22_X1 U2528 ( .A1(n18469), .A2(n18752), .B1(n17830), .B2(n18757), .ZN(
        n3053) );
  OAI22_X1 U2529 ( .A1(n18466), .A2(n18752), .B1(n17831), .B2(n18756), .ZN(
        n3054) );
  OAI22_X1 U2530 ( .A1(n18463), .A2(n18752), .B1(n17832), .B2(n18756), .ZN(
        n3055) );
  OAI22_X1 U2531 ( .A1(n18459), .A2(n18752), .B1(n17833), .B2(n18756), .ZN(
        n3056) );
  OAI22_X1 U2532 ( .A1(n18457), .A2(n18752), .B1(n17834), .B2(n18756), .ZN(
        n3057) );
  OAI22_X1 U2533 ( .A1(n18454), .A2(n18752), .B1(n17835), .B2(n18755), .ZN(
        n3058) );
  OAI22_X1 U2534 ( .A1(n18451), .A2(n18752), .B1(n17836), .B2(n18755), .ZN(
        n3059) );
  OAI22_X1 U2535 ( .A1(n18448), .A2(n18752), .B1(n17837), .B2(n18755), .ZN(
        n3060) );
  OAI22_X1 U2536 ( .A1(n18445), .A2(n18752), .B1(n17838), .B2(n18755), .ZN(
        n3061) );
  OAI22_X1 U2537 ( .A1(n18489), .A2(n18884), .B1(n17942), .B2(n18887), .ZN(
        n3816) );
  OAI22_X1 U2538 ( .A1(n18486), .A2(n18884), .B1(n17943), .B2(n18887), .ZN(
        n3800) );
  OAI22_X1 U2539 ( .A1(n18483), .A2(n18884), .B1(n17944), .B2(n18887), .ZN(
        n3784) );
  OAI22_X1 U2540 ( .A1(n18480), .A2(n18884), .B1(n17945), .B2(n18887), .ZN(
        n3768) );
  OAI22_X1 U2541 ( .A1(n18477), .A2(n18884), .B1(n17946), .B2(n18888), .ZN(
        n3752) );
  OAI22_X1 U2542 ( .A1(n18474), .A2(n18884), .B1(n17947), .B2(n18888), .ZN(
        n3736) );
  OAI22_X1 U2543 ( .A1(n18471), .A2(n18884), .B1(n17948), .B2(n18888), .ZN(
        n3720) );
  OAI22_X1 U2544 ( .A1(n18468), .A2(n18884), .B1(n17949), .B2(n18888), .ZN(
        n3704) );
  OAI22_X1 U2545 ( .A1(n18465), .A2(n18884), .B1(n17950), .B2(n18889), .ZN(
        n3688) );
  OAI22_X1 U2546 ( .A1(n18462), .A2(n18884), .B1(n17951), .B2(n18889), .ZN(
        n3672) );
  OAI22_X1 U2547 ( .A1(n18459), .A2(n18884), .B1(n17952), .B2(n18889), .ZN(
        n3656) );
  OAI22_X1 U2548 ( .A1(n18456), .A2(n18884), .B1(n17953), .B2(n18889), .ZN(
        n3640) );
  OAI22_X1 U2549 ( .A1(n18453), .A2(n18883), .B1(n17954), .B2(n18890), .ZN(
        n3624) );
  OAI22_X1 U2550 ( .A1(n18450), .A2(n18883), .B1(n17955), .B2(n18890), .ZN(
        n3608) );
  OAI22_X1 U2551 ( .A1(n18447), .A2(n18883), .B1(n17956), .B2(n18890), .ZN(
        n3592) );
  OAI22_X1 U2552 ( .A1(n18444), .A2(n18883), .B1(n17957), .B2(n18890), .ZN(
        n3576) );
  OAI22_X1 U2553 ( .A1(n18441), .A2(n18883), .B1(n17958), .B2(n18891), .ZN(
        n3560) );
  OAI22_X1 U2554 ( .A1(n18438), .A2(n18883), .B1(n17959), .B2(n18891), .ZN(
        n3544) );
  OAI22_X1 U2555 ( .A1(n18435), .A2(n18883), .B1(n17960), .B2(n18891), .ZN(
        n3528) );
  OAI22_X1 U2556 ( .A1(n18432), .A2(n18883), .B1(n17961), .B2(n18891), .ZN(
        n3512) );
  OAI22_X1 U2557 ( .A1(n18429), .A2(n18883), .B1(n17962), .B2(n18892), .ZN(
        n3496) );
  OAI22_X1 U2558 ( .A1(n18426), .A2(n18883), .B1(n17963), .B2(n18892), .ZN(
        n3480) );
  OAI22_X1 U2559 ( .A1(n18423), .A2(n18883), .B1(n17964), .B2(n18892), .ZN(
        n3464) );
  OAI22_X1 U2560 ( .A1(n18420), .A2(n18883), .B1(n17965), .B2(n18892), .ZN(
        n3448) );
  OAI22_X1 U2561 ( .A1(n18500), .A2(n18993), .B1(n18031), .B2(n18995), .ZN(
        n8986) );
  OAI22_X1 U2562 ( .A1(n18464), .A2(n18994), .B1(n18043), .B2(n18995), .ZN(
        n8998) );
  OAI22_X1 U2563 ( .A1(n18458), .A2(n18994), .B1(n18045), .B2(n18995), .ZN(
        n9000) );
  OAI22_X1 U2564 ( .A1(n18452), .A2(n18994), .B1(n18047), .B2(n18995), .ZN(
        n9002) );
  OAI22_X1 U2565 ( .A1(n18452), .A2(n18916), .B1(n18063), .B2(n18918), .ZN(
        n3629) );
  OAI22_X1 U2566 ( .A1(n18442), .A2(n18752), .B1(n18203), .B2(n18754), .ZN(
        n3062) );
  OAI22_X1 U2567 ( .A1(n18439), .A2(n18751), .B1(n18204), .B2(n18754), .ZN(
        n3063) );
  OAI22_X1 U2568 ( .A1(n18436), .A2(n18752), .B1(n18205), .B2(n18754), .ZN(
        n3064) );
  OAI22_X1 U2569 ( .A1(n18433), .A2(n18751), .B1(n18206), .B2(n18754), .ZN(
        n3065) );
  OAI22_X1 U2570 ( .A1(n18430), .A2(n18752), .B1(n18207), .B2(n18753), .ZN(
        n3066) );
  OAI22_X1 U2571 ( .A1(n18427), .A2(n18751), .B1(n18208), .B2(n18753), .ZN(
        n3067) );
  OAI22_X1 U2572 ( .A1(n18424), .A2(n18752), .B1(n18209), .B2(n18753), .ZN(
        n3068) );
  OAI22_X1 U2573 ( .A1(n18421), .A2(n18751), .B1(n18210), .B2(n18753), .ZN(
        n3069) );
  OAI22_X1 U2574 ( .A1(n18513), .A2(n18884), .B1(n18243), .B2(n18885), .ZN(
        n3944) );
  OAI22_X1 U2575 ( .A1(n18510), .A2(n18883), .B1(n18244), .B2(n18885), .ZN(
        n3928) );
  OAI22_X1 U2576 ( .A1(n18507), .A2(n18884), .B1(n18245), .B2(n18885), .ZN(
        n3912) );
  OAI22_X1 U2577 ( .A1(n18504), .A2(n18883), .B1(n18246), .B2(n18885), .ZN(
        n3896) );
  OAI22_X1 U2578 ( .A1(n18501), .A2(n18884), .B1(n18247), .B2(n18886), .ZN(
        n3880) );
  OAI22_X1 U2579 ( .A1(n18498), .A2(n18883), .B1(n18248), .B2(n18886), .ZN(
        n3864) );
  OAI22_X1 U2580 ( .A1(n18495), .A2(n18884), .B1(n18249), .B2(n18886), .ZN(
        n3848) );
  OAI22_X1 U2581 ( .A1(n18492), .A2(n18883), .B1(n18250), .B2(n18886), .ZN(
        n3832) );
  OAI22_X1 U2582 ( .A1(n18512), .A2(n19035), .B1(n2494), .B2(n19044), .ZN(
        n9142) );
  OAI22_X1 U2583 ( .A1(n18509), .A2(n19035), .B1(n2485), .B2(n19044), .ZN(
        n9143) );
  OAI22_X1 U2584 ( .A1(n18506), .A2(n19035), .B1(n2476), .B2(n19044), .ZN(
        n9144) );
  OAI22_X1 U2585 ( .A1(n18503), .A2(n19035), .B1(n2467), .B2(n19044), .ZN(
        n9145) );
  OAI22_X1 U2586 ( .A1(n18500), .A2(n19035), .B1(n2458), .B2(n19043), .ZN(
        n9146) );
  OAI22_X1 U2587 ( .A1(n18497), .A2(n19035), .B1(n2449), .B2(n19043), .ZN(
        n9147) );
  OAI22_X1 U2588 ( .A1(n18494), .A2(n19035), .B1(n2440), .B2(n19043), .ZN(
        n9148) );
  OAI22_X1 U2589 ( .A1(n18491), .A2(n19035), .B1(n2431), .B2(n19043), .ZN(
        n9149) );
  OAI22_X1 U2590 ( .A1(n18488), .A2(n19035), .B1(n2422), .B2(n19042), .ZN(
        n9150) );
  OAI22_X1 U2591 ( .A1(n18485), .A2(n19035), .B1(n2413), .B2(n19042), .ZN(
        n9151) );
  OAI22_X1 U2592 ( .A1(n18482), .A2(n19035), .B1(n2404), .B2(n19042), .ZN(
        n9152) );
  OAI22_X1 U2593 ( .A1(n18479), .A2(n19035), .B1(n2395), .B2(n19042), .ZN(
        n9153) );
  OAI22_X1 U2594 ( .A1(n18476), .A2(n19036), .B1(n2386), .B2(n19041), .ZN(
        n9154) );
  OAI22_X1 U2595 ( .A1(n18473), .A2(n19036), .B1(n2377), .B2(n19041), .ZN(
        n9155) );
  OAI22_X1 U2596 ( .A1(n18470), .A2(n19036), .B1(n2368), .B2(n19041), .ZN(
        n9156) );
  OAI22_X1 U2597 ( .A1(n18467), .A2(n19036), .B1(n2359), .B2(n19041), .ZN(
        n9157) );
  OAI22_X1 U2598 ( .A1(n18464), .A2(n19036), .B1(n2350), .B2(n19040), .ZN(
        n9158) );
  OAI22_X1 U2599 ( .A1(n18461), .A2(n19036), .B1(n2341), .B2(n19040), .ZN(
        n9159) );
  OAI22_X1 U2600 ( .A1(n18458), .A2(n19036), .B1(n2332), .B2(n19040), .ZN(
        n9160) );
  OAI22_X1 U2601 ( .A1(n18455), .A2(n19036), .B1(n2323), .B2(n19040), .ZN(
        n9161) );
  OAI22_X1 U2602 ( .A1(n18452), .A2(n19036), .B1(n2314), .B2(n19039), .ZN(
        n9162) );
  OAI22_X1 U2603 ( .A1(n18449), .A2(n19036), .B1(n2305), .B2(n19039), .ZN(
        n9163) );
  OAI22_X1 U2604 ( .A1(n18446), .A2(n19036), .B1(n2296), .B2(n19039), .ZN(
        n9164) );
  OAI22_X1 U2605 ( .A1(n18443), .A2(n19036), .B1(n2287), .B2(n19039), .ZN(
        n9165) );
  OAI22_X1 U2606 ( .A1(n18440), .A2(n19035), .B1(n2278), .B2(n19038), .ZN(
        n9166) );
  OAI22_X1 U2607 ( .A1(n18437), .A2(n19036), .B1(n2269), .B2(n19038), .ZN(
        n9167) );
  OAI22_X1 U2608 ( .A1(n18434), .A2(n19035), .B1(n2260), .B2(n19038), .ZN(
        n9168) );
  OAI22_X1 U2609 ( .A1(n18431), .A2(n19036), .B1(n2251), .B2(n19038), .ZN(
        n9169) );
  OAI22_X1 U2610 ( .A1(n18428), .A2(n19035), .B1(n2242), .B2(n19037), .ZN(
        n9170) );
  OAI22_X1 U2611 ( .A1(n18425), .A2(n19036), .B1(n2233), .B2(n19037), .ZN(
        n9171) );
  OAI22_X1 U2612 ( .A1(n18422), .A2(n19035), .B1(n2224), .B2(n19037), .ZN(
        n9172) );
  OAI22_X1 U2613 ( .A1(n18419), .A2(n19036), .B1(n2215), .B2(n19037), .ZN(
        n9173) );
  OAI22_X1 U2614 ( .A1(n18483), .A2(n18861), .B1(n17966), .B2(n18865), .ZN(
        n3368) );
  OAI22_X1 U2615 ( .A1(n18480), .A2(n18861), .B1(n17967), .B2(n18865), .ZN(
        n3369) );
  OAI22_X1 U2616 ( .A1(n18477), .A2(n18862), .B1(n17968), .B2(n18865), .ZN(
        n3370) );
  OAI22_X1 U2617 ( .A1(n18474), .A2(n18862), .B1(n17969), .B2(n18864), .ZN(
        n3371) );
  OAI22_X1 U2618 ( .A1(n18471), .A2(n18862), .B1(n17970), .B2(n18865), .ZN(
        n3372) );
  OAI22_X1 U2619 ( .A1(n18468), .A2(n18862), .B1(n17971), .B2(n18866), .ZN(
        n3373) );
  OAI22_X1 U2620 ( .A1(n18465), .A2(n18862), .B1(n17972), .B2(n18866), .ZN(
        n3374) );
  OAI22_X1 U2621 ( .A1(n18462), .A2(n18862), .B1(n17973), .B2(n18864), .ZN(
        n3375) );
  OAI22_X1 U2622 ( .A1(n18459), .A2(n18862), .B1(n17974), .B2(n18863), .ZN(
        n3376) );
  OAI22_X1 U2623 ( .A1(n18456), .A2(n18862), .B1(n17975), .B2(n18863), .ZN(
        n3377) );
  OAI22_X1 U2624 ( .A1(n18453), .A2(n18862), .B1(n17976), .B2(n18864), .ZN(
        n3378) );
  OAI22_X1 U2625 ( .A1(n18450), .A2(n18862), .B1(n17977), .B2(n18864), .ZN(
        n3379) );
  OAI22_X1 U2626 ( .A1(n18447), .A2(n18862), .B1(n17978), .B2(n18863), .ZN(
        n3380) );
  OAI22_X1 U2627 ( .A1(n18444), .A2(n18862), .B1(n17979), .B2(n18863), .ZN(
        n3381) );
  OAI22_X1 U2628 ( .A1(n18513), .A2(n18795), .B1(n18171), .B2(n18804), .ZN(
        n3166) );
  OAI22_X1 U2629 ( .A1(n18510), .A2(n18795), .B1(n18172), .B2(n18804), .ZN(
        n3167) );
  OAI22_X1 U2630 ( .A1(n18507), .A2(n18795), .B1(n18173), .B2(n18804), .ZN(
        n3168) );
  OAI22_X1 U2631 ( .A1(n18504), .A2(n18795), .B1(n18174), .B2(n18804), .ZN(
        n3169) );
  OAI22_X1 U2632 ( .A1(n18501), .A2(n18795), .B1(n18175), .B2(n18803), .ZN(
        n3170) );
  OAI22_X1 U2633 ( .A1(n18498), .A2(n18795), .B1(n18176), .B2(n18803), .ZN(
        n3171) );
  OAI22_X1 U2634 ( .A1(n18492), .A2(n18795), .B1(n18178), .B2(n18803), .ZN(
        n3173) );
  OAI22_X1 U2635 ( .A1(n18489), .A2(n18795), .B1(n18179), .B2(n18802), .ZN(
        n3174) );
  OAI22_X1 U2636 ( .A1(n18486), .A2(n18795), .B1(n18180), .B2(n18802), .ZN(
        n3175) );
  OAI22_X1 U2637 ( .A1(n18483), .A2(n18795), .B1(n18181), .B2(n18802), .ZN(
        n3176) );
  OAI22_X1 U2638 ( .A1(n18480), .A2(n18795), .B1(n18182), .B2(n18802), .ZN(
        n3177) );
  OAI22_X1 U2639 ( .A1(n18477), .A2(n18796), .B1(n18183), .B2(n18801), .ZN(
        n3178) );
  OAI22_X1 U2640 ( .A1(n18474), .A2(n18796), .B1(n18184), .B2(n18801), .ZN(
        n3179) );
  OAI22_X1 U2641 ( .A1(n18471), .A2(n18796), .B1(n18185), .B2(n18801), .ZN(
        n3180) );
  OAI22_X1 U2642 ( .A1(n18468), .A2(n18796), .B1(n18186), .B2(n18801), .ZN(
        n3181) );
  OAI22_X1 U2643 ( .A1(n18465), .A2(n18796), .B1(n18187), .B2(n18800), .ZN(
        n3182) );
  OAI22_X1 U2644 ( .A1(n18462), .A2(n18796), .B1(n18188), .B2(n18800), .ZN(
        n3183) );
  OAI22_X1 U2645 ( .A1(n18459), .A2(n18796), .B1(n18189), .B2(n18800), .ZN(
        n3184) );
  OAI22_X1 U2646 ( .A1(n18456), .A2(n18796), .B1(n18190), .B2(n18800), .ZN(
        n3185) );
  OAI22_X1 U2647 ( .A1(n18453), .A2(n18796), .B1(n18191), .B2(n18799), .ZN(
        n3186) );
  OAI22_X1 U2648 ( .A1(n18450), .A2(n18796), .B1(n18192), .B2(n18799), .ZN(
        n3187) );
  OAI22_X1 U2649 ( .A1(n18447), .A2(n18796), .B1(n18193), .B2(n18799), .ZN(
        n3188) );
  OAI22_X1 U2650 ( .A1(n18444), .A2(n18796), .B1(n18194), .B2(n18799), .ZN(
        n3189) );
  OAI22_X1 U2651 ( .A1(n18441), .A2(n18795), .B1(n18315), .B2(n18798), .ZN(
        n3190) );
  OAI22_X1 U2652 ( .A1(n18438), .A2(n18796), .B1(n18316), .B2(n18798), .ZN(
        n3191) );
  OAI22_X1 U2653 ( .A1(n18435), .A2(n18795), .B1(n18317), .B2(n18798), .ZN(
        n3192) );
  OAI22_X1 U2654 ( .A1(n18432), .A2(n18796), .B1(n18318), .B2(n18798), .ZN(
        n3193) );
  OAI22_X1 U2655 ( .A1(n18429), .A2(n18795), .B1(n18319), .B2(n18797), .ZN(
        n3194) );
  OAI22_X1 U2656 ( .A1(n18426), .A2(n18796), .B1(n18320), .B2(n18797), .ZN(
        n3195) );
  OAI22_X1 U2657 ( .A1(n18423), .A2(n18795), .B1(n18321), .B2(n18797), .ZN(
        n3196) );
  OAI22_X1 U2658 ( .A1(n18420), .A2(n18796), .B1(n18322), .B2(n18797), .ZN(
        n3197) );
  OAI22_X1 U2659 ( .A1(n18495), .A2(n18806), .B1(n17877), .B2(n18814), .ZN(
        n3204) );
  OAI22_X1 U2660 ( .A1(n18495), .A2(n18795), .B1(n18177), .B2(n18803), .ZN(
        n3172) );
  OAI22_X1 U2661 ( .A1(n18490), .A2(n18719), .B1(n2427), .B2(n18720), .ZN(
        n2908) );
  OAI22_X1 U2662 ( .A1(n18487), .A2(n18718), .B1(n2418), .B2(n18720), .ZN(
        n2907) );
  OAI22_X1 U2663 ( .A1(n18484), .A2(n18719), .B1(n2409), .B2(n18720), .ZN(
        n2906) );
  OAI22_X1 U2664 ( .A1(n18481), .A2(n18718), .B1(n2400), .B2(n18720), .ZN(
        n2905) );
  OAI22_X1 U2665 ( .A1(n18478), .A2(n18719), .B1(n2391), .B2(n18721), .ZN(
        n2904) );
  OAI22_X1 U2666 ( .A1(n18475), .A2(n18718), .B1(n2382), .B2(n18721), .ZN(
        n2903) );
  OAI22_X1 U2667 ( .A1(n18472), .A2(n18719), .B1(n2373), .B2(n18721), .ZN(
        n2902) );
  OAI22_X1 U2668 ( .A1(n18469), .A2(n18718), .B1(n2364), .B2(n18721), .ZN(
        n2901) );
  OAI22_X1 U2669 ( .A1(n18466), .A2(n18719), .B1(n2355), .B2(n18722), .ZN(
        n2900) );
  OAI22_X1 U2670 ( .A1(n18463), .A2(n18719), .B1(n2346), .B2(n18722), .ZN(
        n2899) );
  OAI22_X1 U2671 ( .A1(n18460), .A2(n18719), .B1(n2337), .B2(n18722), .ZN(
        n2898) );
  OAI22_X1 U2672 ( .A1(n18457), .A2(n18719), .B1(n2328), .B2(n18722), .ZN(
        n2897) );
  OAI22_X1 U2673 ( .A1(n18454), .A2(n18719), .B1(n2319), .B2(n18723), .ZN(
        n2896) );
  OAI22_X1 U2674 ( .A1(n18451), .A2(n18719), .B1(n2310), .B2(n18723), .ZN(
        n2895) );
  OAI22_X1 U2675 ( .A1(n18448), .A2(n18719), .B1(n2301), .B2(n18723), .ZN(
        n2894) );
  OAI22_X1 U2676 ( .A1(n18445), .A2(n18719), .B1(n2292), .B2(n18723), .ZN(
        n2893) );
  OAI22_X1 U2677 ( .A1(n18442), .A2(n18719), .B1(n2283), .B2(n18724), .ZN(
        n2892) );
  OAI22_X1 U2678 ( .A1(n18439), .A2(n18719), .B1(n2274), .B2(n18724), .ZN(
        n2891) );
  OAI22_X1 U2679 ( .A1(n18436), .A2(n18719), .B1(n2265), .B2(n18724), .ZN(
        n2890) );
  OAI22_X1 U2680 ( .A1(n18433), .A2(n18719), .B1(n2256), .B2(n18724), .ZN(
        n2889) );
  OAI22_X1 U2681 ( .A1(n18430), .A2(n18718), .B1(n2247), .B2(n18725), .ZN(
        n2888) );
  OAI22_X1 U2682 ( .A1(n18427), .A2(n18718), .B1(n2238), .B2(n18725), .ZN(
        n2887) );
  OAI22_X1 U2683 ( .A1(n18424), .A2(n18718), .B1(n2229), .B2(n18725), .ZN(
        n2886) );
  OAI22_X1 U2684 ( .A1(n18421), .A2(n18718), .B1(n2220), .B2(n18725), .ZN(
        n2885) );
  OAI22_X1 U2685 ( .A1(n18514), .A2(n18718), .B1(n2499), .B2(n18726), .ZN(
        n2884) );
  OAI22_X1 U2686 ( .A1(n18511), .A2(n18718), .B1(n2490), .B2(n18726), .ZN(
        n2883) );
  OAI22_X1 U2687 ( .A1(n18508), .A2(n18718), .B1(n2481), .B2(n18726), .ZN(
        n2882) );
  OAI22_X1 U2688 ( .A1(n18505), .A2(n18718), .B1(n2472), .B2(n18726), .ZN(
        n2881) );
  OAI22_X1 U2689 ( .A1(n18502), .A2(n18718), .B1(n2463), .B2(n18727), .ZN(
        n2880) );
  OAI22_X1 U2690 ( .A1(n18499), .A2(n18718), .B1(n2454), .B2(n18727), .ZN(
        n2879) );
  OAI22_X1 U2691 ( .A1(n18496), .A2(n18718), .B1(n2445), .B2(n18727), .ZN(
        n2878) );
  OAI22_X1 U2692 ( .A1(n18493), .A2(n18718), .B1(n2436), .B2(n18727), .ZN(
        n2877) );
  OAI22_X1 U2693 ( .A1(n18488), .A2(n18928), .B1(n2423), .B2(n18931), .ZN(
        n3824) );
  OAI22_X1 U2694 ( .A1(n18485), .A2(n18928), .B1(n2414), .B2(n18931), .ZN(
        n3808) );
  OAI22_X1 U2695 ( .A1(n18482), .A2(n18928), .B1(n2405), .B2(n18931), .ZN(
        n3792) );
  OAI22_X1 U2696 ( .A1(n18479), .A2(n18928), .B1(n2396), .B2(n18931), .ZN(
        n3776) );
  OAI22_X1 U2697 ( .A1(n18476), .A2(n18928), .B1(n2387), .B2(n18932), .ZN(
        n3760) );
  OAI22_X1 U2698 ( .A1(n18473), .A2(n18928), .B1(n2378), .B2(n18932), .ZN(
        n3744) );
  OAI22_X1 U2699 ( .A1(n18470), .A2(n18928), .B1(n2369), .B2(n18932), .ZN(
        n3728) );
  OAI22_X1 U2700 ( .A1(n18467), .A2(n18928), .B1(n2360), .B2(n18932), .ZN(
        n3712) );
  OAI22_X1 U2701 ( .A1(n18464), .A2(n18928), .B1(n2351), .B2(n18933), .ZN(
        n3696) );
  OAI22_X1 U2702 ( .A1(n18461), .A2(n18928), .B1(n2342), .B2(n18933), .ZN(
        n3680) );
  OAI22_X1 U2703 ( .A1(n18458), .A2(n18928), .B1(n2333), .B2(n18933), .ZN(
        n3664) );
  OAI22_X1 U2704 ( .A1(n18455), .A2(n18928), .B1(n2324), .B2(n18933), .ZN(
        n3648) );
  OAI22_X1 U2705 ( .A1(n18452), .A2(n18927), .B1(n2315), .B2(n18934), .ZN(
        n3632) );
  OAI22_X1 U2706 ( .A1(n18449), .A2(n18927), .B1(n2306), .B2(n18934), .ZN(
        n3616) );
  OAI22_X1 U2707 ( .A1(n18446), .A2(n18927), .B1(n2297), .B2(n18934), .ZN(
        n3600) );
  OAI22_X1 U2708 ( .A1(n18443), .A2(n18927), .B1(n2288), .B2(n18934), .ZN(
        n3584) );
  OAI22_X1 U2709 ( .A1(n18440), .A2(n18927), .B1(n2279), .B2(n18935), .ZN(
        n3568) );
  OAI22_X1 U2710 ( .A1(n18437), .A2(n18927), .B1(n2270), .B2(n18935), .ZN(
        n3552) );
  OAI22_X1 U2711 ( .A1(n18434), .A2(n18927), .B1(n2261), .B2(n18935), .ZN(
        n3536) );
  OAI22_X1 U2712 ( .A1(n18431), .A2(n18927), .B1(n2252), .B2(n18935), .ZN(
        n3520) );
  OAI22_X1 U2713 ( .A1(n18428), .A2(n18927), .B1(n2243), .B2(n18936), .ZN(
        n3504) );
  OAI22_X1 U2714 ( .A1(n18425), .A2(n18927), .B1(n2234), .B2(n18936), .ZN(
        n3488) );
  OAI22_X1 U2715 ( .A1(n18422), .A2(n18927), .B1(n2225), .B2(n18936), .ZN(
        n3472) );
  OAI22_X1 U2716 ( .A1(n18419), .A2(n18927), .B1(n2216), .B2(n18936), .ZN(
        n3456) );
  OAI22_X1 U2717 ( .A1(n18489), .A2(n18895), .B1(n2428), .B2(n18898), .ZN(
        n3818) );
  OAI22_X1 U2718 ( .A1(n18486), .A2(n18895), .B1(n2419), .B2(n18898), .ZN(
        n3802) );
  OAI22_X1 U2719 ( .A1(n18483), .A2(n18895), .B1(n2410), .B2(n18898), .ZN(
        n3786) );
  OAI22_X1 U2720 ( .A1(n18480), .A2(n18895), .B1(n2401), .B2(n18898), .ZN(
        n3770) );
  OAI22_X1 U2721 ( .A1(n18477), .A2(n18895), .B1(n2392), .B2(n18899), .ZN(
        n3754) );
  OAI22_X1 U2722 ( .A1(n18474), .A2(n18895), .B1(n2383), .B2(n18899), .ZN(
        n3738) );
  OAI22_X1 U2723 ( .A1(n18471), .A2(n18895), .B1(n2374), .B2(n18899), .ZN(
        n3722) );
  OAI22_X1 U2724 ( .A1(n18468), .A2(n18895), .B1(n2365), .B2(n18899), .ZN(
        n3706) );
  OAI22_X1 U2725 ( .A1(n18465), .A2(n18895), .B1(n2356), .B2(n18900), .ZN(
        n3690) );
  OAI22_X1 U2726 ( .A1(n18462), .A2(n18895), .B1(n2347), .B2(n18900), .ZN(
        n3674) );
  OAI22_X1 U2727 ( .A1(n18458), .A2(n18895), .B1(n2338), .B2(n18900), .ZN(
        n3658) );
  OAI22_X1 U2728 ( .A1(n18456), .A2(n18895), .B1(n2329), .B2(n18900), .ZN(
        n3642) );
  OAI22_X1 U2729 ( .A1(n18453), .A2(n18894), .B1(n2320), .B2(n18901), .ZN(
        n3626) );
  OAI22_X1 U2730 ( .A1(n18450), .A2(n18894), .B1(n2311), .B2(n18901), .ZN(
        n3610) );
  OAI22_X1 U2731 ( .A1(n18447), .A2(n18894), .B1(n2302), .B2(n18901), .ZN(
        n3594) );
  OAI22_X1 U2732 ( .A1(n18444), .A2(n18894), .B1(n2293), .B2(n18901), .ZN(
        n3578) );
  OAI22_X1 U2733 ( .A1(n18441), .A2(n18894), .B1(n2284), .B2(n18902), .ZN(
        n3562) );
  OAI22_X1 U2734 ( .A1(n18438), .A2(n18894), .B1(n2275), .B2(n18902), .ZN(
        n3546) );
  OAI22_X1 U2735 ( .A1(n18435), .A2(n18894), .B1(n2266), .B2(n18902), .ZN(
        n3530) );
  OAI22_X1 U2736 ( .A1(n18432), .A2(n18894), .B1(n2257), .B2(n18902), .ZN(
        n3514) );
  OAI22_X1 U2737 ( .A1(n18429), .A2(n18894), .B1(n2248), .B2(n18903), .ZN(
        n3498) );
  OAI22_X1 U2738 ( .A1(n18426), .A2(n18894), .B1(n2239), .B2(n18903), .ZN(
        n3482) );
  OAI22_X1 U2739 ( .A1(n18423), .A2(n18894), .B1(n2230), .B2(n18903), .ZN(
        n3466) );
  OAI22_X1 U2740 ( .A1(n18420), .A2(n18894), .B1(n2221), .B2(n18903), .ZN(
        n3450) );
  OAI22_X1 U2741 ( .A1(n18512), .A2(n18928), .B1(n2495), .B2(n18929), .ZN(
        n3952) );
  OAI22_X1 U2742 ( .A1(n18509), .A2(n18927), .B1(n2486), .B2(n18929), .ZN(
        n3936) );
  OAI22_X1 U2743 ( .A1(n18506), .A2(n18928), .B1(n2477), .B2(n18929), .ZN(
        n3920) );
  OAI22_X1 U2744 ( .A1(n18503), .A2(n18927), .B1(n2468), .B2(n18929), .ZN(
        n3904) );
  OAI22_X1 U2745 ( .A1(n18500), .A2(n18928), .B1(n2459), .B2(n18930), .ZN(
        n3888) );
  OAI22_X1 U2746 ( .A1(n18497), .A2(n18927), .B1(n2450), .B2(n18930), .ZN(
        n3872) );
  OAI22_X1 U2747 ( .A1(n18494), .A2(n18928), .B1(n2441), .B2(n18930), .ZN(
        n3856) );
  OAI22_X1 U2748 ( .A1(n18491), .A2(n18927), .B1(n2432), .B2(n18930), .ZN(
        n3840) );
  OAI22_X1 U2749 ( .A1(n18513), .A2(n18895), .B1(n2500), .B2(n18896), .ZN(
        n3946) );
  OAI22_X1 U2750 ( .A1(n18510), .A2(n18894), .B1(n2491), .B2(n18896), .ZN(
        n3930) );
  OAI22_X1 U2751 ( .A1(n18507), .A2(n18895), .B1(n2482), .B2(n18896), .ZN(
        n3914) );
  OAI22_X1 U2752 ( .A1(n18504), .A2(n18894), .B1(n2473), .B2(n18896), .ZN(
        n3898) );
  OAI22_X1 U2753 ( .A1(n18501), .A2(n18895), .B1(n2464), .B2(n18897), .ZN(
        n3882) );
  OAI22_X1 U2754 ( .A1(n18498), .A2(n18894), .B1(n2455), .B2(n18897), .ZN(
        n3866) );
  OAI22_X1 U2755 ( .A1(n18495), .A2(n18895), .B1(n2446), .B2(n18897), .ZN(
        n3850) );
  OAI22_X1 U2756 ( .A1(n18492), .A2(n18894), .B1(n2437), .B2(n18897), .ZN(
        n3834) );
  OAI22_X1 U2757 ( .A1(n18514), .A2(n18729), .B1(n2498), .B2(n18738), .ZN(
        n2942) );
  OAI22_X1 U2758 ( .A1(n18511), .A2(n18729), .B1(n2489), .B2(n18738), .ZN(
        n2943) );
  OAI22_X1 U2759 ( .A1(n18508), .A2(n18729), .B1(n2480), .B2(n18738), .ZN(
        n2944) );
  OAI22_X1 U2760 ( .A1(n18505), .A2(n18729), .B1(n2471), .B2(n18737), .ZN(
        n2945) );
  OAI22_X1 U2761 ( .A1(n18502), .A2(n18729), .B1(n2462), .B2(n18737), .ZN(
        n2946) );
  OAI22_X1 U2762 ( .A1(n18499), .A2(n18729), .B1(n2453), .B2(n18737), .ZN(
        n2947) );
  OAI22_X1 U2763 ( .A1(n18496), .A2(n18729), .B1(n2444), .B2(n18737), .ZN(
        n2948) );
  OAI22_X1 U2764 ( .A1(n18493), .A2(n18729), .B1(n2435), .B2(n18736), .ZN(
        n2949) );
  OAI22_X1 U2765 ( .A1(n18490), .A2(n18729), .B1(n2426), .B2(n18736), .ZN(
        n2950) );
  OAI22_X1 U2766 ( .A1(n18487), .A2(n18729), .B1(n2417), .B2(n18736), .ZN(
        n2951) );
  OAI22_X1 U2767 ( .A1(n18484), .A2(n18729), .B1(n2408), .B2(n18736), .ZN(
        n2952) );
  OAI22_X1 U2768 ( .A1(n18481), .A2(n18730), .B1(n2399), .B2(n18735), .ZN(
        n2953) );
  OAI22_X1 U2769 ( .A1(n18478), .A2(n18730), .B1(n2390), .B2(n18735), .ZN(
        n2954) );
  OAI22_X1 U2770 ( .A1(n18475), .A2(n18730), .B1(n2381), .B2(n18735), .ZN(
        n2955) );
  OAI22_X1 U2771 ( .A1(n18472), .A2(n18730), .B1(n2372), .B2(n18735), .ZN(
        n2956) );
  OAI22_X1 U2772 ( .A1(n18469), .A2(n18730), .B1(n2363), .B2(n18734), .ZN(
        n2957) );
  OAI22_X1 U2773 ( .A1(n18466), .A2(n18730), .B1(n2354), .B2(n18734), .ZN(
        n2958) );
  OAI22_X1 U2774 ( .A1(n18463), .A2(n18730), .B1(n2345), .B2(n18734), .ZN(
        n2959) );
  OAI22_X1 U2775 ( .A1(n18460), .A2(n18730), .B1(n2336), .B2(n18734), .ZN(
        n2960) );
  OAI22_X1 U2776 ( .A1(n18457), .A2(n18730), .B1(n2327), .B2(n18733), .ZN(
        n2961) );
  OAI22_X1 U2777 ( .A1(n18454), .A2(n18729), .B1(n2318), .B2(n18738), .ZN(
        n18386) );
  OAI22_X1 U2778 ( .A1(n18451), .A2(n18730), .B1(n2309), .B2(n18733), .ZN(
        n2963) );
  OAI22_X1 U2779 ( .A1(n18448), .A2(n18730), .B1(n2300), .B2(n18733), .ZN(
        n2964) );
  OAI22_X1 U2780 ( .A1(n18445), .A2(n18730), .B1(n2291), .B2(n18733), .ZN(
        n2965) );
  OAI22_X1 U2781 ( .A1(n18488), .A2(n18906), .B1(n2429), .B2(n18909), .ZN(
        n3820) );
  OAI22_X1 U2782 ( .A1(n18485), .A2(n18906), .B1(n2420), .B2(n18909), .ZN(
        n3804) );
  OAI22_X1 U2783 ( .A1(n18482), .A2(n18906), .B1(n2411), .B2(n18909), .ZN(
        n3788) );
  OAI22_X1 U2784 ( .A1(n18479), .A2(n18906), .B1(n2402), .B2(n18909), .ZN(
        n3772) );
  OAI22_X1 U2785 ( .A1(n18476), .A2(n18906), .B1(n2393), .B2(n18910), .ZN(
        n3756) );
  OAI22_X1 U2786 ( .A1(n18473), .A2(n18906), .B1(n2384), .B2(n18910), .ZN(
        n3740) );
  OAI22_X1 U2787 ( .A1(n18470), .A2(n18906), .B1(n2375), .B2(n18910), .ZN(
        n3724) );
  OAI22_X1 U2788 ( .A1(n18467), .A2(n18906), .B1(n2366), .B2(n18910), .ZN(
        n3708) );
  OAI22_X1 U2789 ( .A1(n18464), .A2(n18906), .B1(n2357), .B2(n18911), .ZN(
        n3692) );
  OAI22_X1 U2790 ( .A1(n18461), .A2(n18906), .B1(n2348), .B2(n18911), .ZN(
        n3676) );
  OAI22_X1 U2791 ( .A1(n18460), .A2(n18905), .B1(n2339), .B2(n18914), .ZN(
        n18387) );
  OAI22_X1 U2792 ( .A1(n18455), .A2(n18906), .B1(n2330), .B2(n18911), .ZN(
        n3644) );
  OAI22_X1 U2793 ( .A1(n18452), .A2(n18906), .B1(n2321), .B2(n18911), .ZN(
        n3628) );
  OAI22_X1 U2794 ( .A1(n18449), .A2(n18905), .B1(n2312), .B2(n18912), .ZN(
        n3612) );
  OAI22_X1 U2795 ( .A1(n18446), .A2(n18905), .B1(n2303), .B2(n18912), .ZN(
        n3596) );
  OAI22_X1 U2796 ( .A1(n18443), .A2(n18905), .B1(n2294), .B2(n18912), .ZN(
        n3580) );
  OAI22_X1 U2797 ( .A1(n18440), .A2(n18905), .B1(n2285), .B2(n18912), .ZN(
        n3564) );
  OAI22_X1 U2798 ( .A1(n18437), .A2(n18905), .B1(n2276), .B2(n18913), .ZN(
        n3548) );
  OAI22_X1 U2799 ( .A1(n18434), .A2(n18905), .B1(n2267), .B2(n18913), .ZN(
        n3532) );
  OAI22_X1 U2800 ( .A1(n18431), .A2(n18905), .B1(n2258), .B2(n18913), .ZN(
        n3516) );
  OAI22_X1 U2801 ( .A1(n18428), .A2(n18905), .B1(n2249), .B2(n18913), .ZN(
        n3500) );
  OAI22_X1 U2802 ( .A1(n18425), .A2(n18905), .B1(n2240), .B2(n18914), .ZN(
        n3484) );
  OAI22_X1 U2803 ( .A1(n18422), .A2(n18905), .B1(n2231), .B2(n18914), .ZN(
        n3468) );
  OAI22_X1 U2804 ( .A1(n18419), .A2(n18905), .B1(n2222), .B2(n18914), .ZN(
        n3452) );
  OAI22_X1 U2805 ( .A1(n18514), .A2(n18740), .B1(n2497), .B2(n18749), .ZN(
        n2974) );
  OAI22_X1 U2806 ( .A1(n18511), .A2(n18740), .B1(n2488), .B2(n18749), .ZN(
        n2975) );
  OAI22_X1 U2807 ( .A1(n18508), .A2(n18740), .B1(n2479), .B2(n18749), .ZN(
        n2976) );
  OAI22_X1 U2808 ( .A1(n18505), .A2(n18740), .B1(n2470), .B2(n18749), .ZN(
        n2977) );
  OAI22_X1 U2809 ( .A1(n18502), .A2(n18740), .B1(n2461), .B2(n18748), .ZN(
        n2978) );
  OAI22_X1 U2810 ( .A1(n18499), .A2(n18740), .B1(n2452), .B2(n18748), .ZN(
        n2979) );
  OAI22_X1 U2811 ( .A1(n18496), .A2(n18740), .B1(n2443), .B2(n18748), .ZN(
        n2980) );
  OAI22_X1 U2812 ( .A1(n18493), .A2(n18740), .B1(n2434), .B2(n18748), .ZN(
        n2981) );
  OAI22_X1 U2813 ( .A1(n18490), .A2(n18740), .B1(n2425), .B2(n18747), .ZN(
        n2982) );
  OAI22_X1 U2814 ( .A1(n18487), .A2(n18740), .B1(n2416), .B2(n18747), .ZN(
        n2983) );
  OAI22_X1 U2815 ( .A1(n18484), .A2(n18740), .B1(n2407), .B2(n18747), .ZN(
        n2984) );
  OAI22_X1 U2816 ( .A1(n18481), .A2(n18740), .B1(n2398), .B2(n18747), .ZN(
        n2985) );
  OAI22_X1 U2817 ( .A1(n18478), .A2(n18741), .B1(n2389), .B2(n18746), .ZN(
        n2986) );
  OAI22_X1 U2818 ( .A1(n18475), .A2(n18741), .B1(n2380), .B2(n18746), .ZN(
        n2987) );
  OAI22_X1 U2819 ( .A1(n18472), .A2(n18741), .B1(n2371), .B2(n18746), .ZN(
        n2988) );
  OAI22_X1 U2820 ( .A1(n18469), .A2(n18741), .B1(n2362), .B2(n18746), .ZN(
        n2989) );
  OAI22_X1 U2821 ( .A1(n18466), .A2(n18741), .B1(n2353), .B2(n18745), .ZN(
        n2990) );
  OAI22_X1 U2822 ( .A1(n18463), .A2(n18741), .B1(n2344), .B2(n18745), .ZN(
        n2991) );
  OAI22_X1 U2823 ( .A1(n18460), .A2(n18741), .B1(n2335), .B2(n18745), .ZN(
        n2992) );
  OAI22_X1 U2824 ( .A1(n18457), .A2(n18741), .B1(n2326), .B2(n18745), .ZN(
        n2993) );
  OAI22_X1 U2825 ( .A1(n18454), .A2(n18741), .B1(n2317), .B2(n18744), .ZN(
        n2994) );
  OAI22_X1 U2826 ( .A1(n18451), .A2(n18741), .B1(n2308), .B2(n18744), .ZN(
        n2995) );
  OAI22_X1 U2827 ( .A1(n18448), .A2(n18741), .B1(n2299), .B2(n18744), .ZN(
        n2996) );
  OAI22_X1 U2828 ( .A1(n18445), .A2(n18741), .B1(n2290), .B2(n18744), .ZN(
        n2997) );
  OAI22_X1 U2829 ( .A1(n18512), .A2(n19015), .B1(n2502), .B2(n19024), .ZN(
        n9046) );
  OAI22_X1 U2830 ( .A1(n18509), .A2(n19015), .B1(n2493), .B2(n19024), .ZN(
        n9047) );
  OAI22_X1 U2831 ( .A1(n18506), .A2(n19015), .B1(n2484), .B2(n19024), .ZN(
        n9048) );
  OAI22_X1 U2832 ( .A1(n18503), .A2(n19015), .B1(n2475), .B2(n19024), .ZN(
        n9049) );
  OAI22_X1 U2833 ( .A1(n18500), .A2(n19015), .B1(n2466), .B2(n19023), .ZN(
        n9050) );
  OAI22_X1 U2834 ( .A1(n18497), .A2(n19015), .B1(n2457), .B2(n19023), .ZN(
        n9051) );
  OAI22_X1 U2835 ( .A1(n18494), .A2(n19015), .B1(n2448), .B2(n19023), .ZN(
        n9052) );
  OAI22_X1 U2836 ( .A1(n18491), .A2(n19015), .B1(n2439), .B2(n19023), .ZN(
        n9053) );
  OAI22_X1 U2837 ( .A1(n18488), .A2(n19015), .B1(n2430), .B2(n19022), .ZN(
        n9054) );
  OAI22_X1 U2838 ( .A1(n18485), .A2(n19015), .B1(n2421), .B2(n19022), .ZN(
        n9055) );
  OAI22_X1 U2839 ( .A1(n18482), .A2(n19015), .B1(n2412), .B2(n19022), .ZN(
        n9056) );
  OAI22_X1 U2840 ( .A1(n18479), .A2(n19015), .B1(n2403), .B2(n19022), .ZN(
        n9057) );
  OAI22_X1 U2841 ( .A1(n18476), .A2(n19016), .B1(n2394), .B2(n19021), .ZN(
        n9058) );
  OAI22_X1 U2842 ( .A1(n18473), .A2(n19016), .B1(n2385), .B2(n19021), .ZN(
        n9059) );
  OAI22_X1 U2843 ( .A1(n18470), .A2(n19016), .B1(n2376), .B2(n19021), .ZN(
        n9060) );
  OAI22_X1 U2844 ( .A1(n18467), .A2(n19016), .B1(n2367), .B2(n19021), .ZN(
        n9061) );
  OAI22_X1 U2845 ( .A1(n18464), .A2(n19016), .B1(n2358), .B2(n19020), .ZN(
        n9062) );
  OAI22_X1 U2846 ( .A1(n18461), .A2(n19016), .B1(n2349), .B2(n19020), .ZN(
        n9063) );
  OAI22_X1 U2847 ( .A1(n18458), .A2(n19016), .B1(n2340), .B2(n19020), .ZN(
        n9064) );
  OAI22_X1 U2848 ( .A1(n18455), .A2(n19016), .B1(n2331), .B2(n19020), .ZN(
        n9065) );
  OAI22_X1 U2849 ( .A1(n18452), .A2(n19016), .B1(n2322), .B2(n19019), .ZN(
        n9066) );
  OAI22_X1 U2850 ( .A1(n18449), .A2(n19016), .B1(n2313), .B2(n19019), .ZN(
        n9067) );
  OAI22_X1 U2851 ( .A1(n18446), .A2(n19016), .B1(n2304), .B2(n19019), .ZN(
        n9068) );
  OAI22_X1 U2852 ( .A1(n18443), .A2(n19016), .B1(n2295), .B2(n19019), .ZN(
        n9069) );
  OAI22_X1 U2853 ( .A1(n18442), .A2(n18729), .B1(n2282), .B2(n18732), .ZN(
        n2966) );
  OAI22_X1 U2854 ( .A1(n18439), .A2(n18730), .B1(n2273), .B2(n18732), .ZN(
        n2967) );
  OAI22_X1 U2855 ( .A1(n18436), .A2(n18729), .B1(n2264), .B2(n18732), .ZN(
        n2968) );
  OAI22_X1 U2856 ( .A1(n18433), .A2(n18730), .B1(n2255), .B2(n18732), .ZN(
        n2969) );
  OAI22_X1 U2857 ( .A1(n18430), .A2(n18729), .B1(n2246), .B2(n18731), .ZN(
        n2970) );
  OAI22_X1 U2858 ( .A1(n18427), .A2(n18730), .B1(n2237), .B2(n18731), .ZN(
        n2971) );
  OAI22_X1 U2859 ( .A1(n18424), .A2(n18729), .B1(n2228), .B2(n18731), .ZN(
        n2972) );
  OAI22_X1 U2860 ( .A1(n18421), .A2(n18730), .B1(n2219), .B2(n18731), .ZN(
        n2973) );
  OAI22_X1 U2861 ( .A1(n18512), .A2(n18906), .B1(n2501), .B2(n18907), .ZN(
        n3948) );
  OAI22_X1 U2862 ( .A1(n18509), .A2(n18905), .B1(n2492), .B2(n18907), .ZN(
        n3932) );
  OAI22_X1 U2863 ( .A1(n18506), .A2(n18906), .B1(n2483), .B2(n18907), .ZN(
        n3916) );
  OAI22_X1 U2864 ( .A1(n18503), .A2(n18905), .B1(n2474), .B2(n18907), .ZN(
        n3900) );
  OAI22_X1 U2865 ( .A1(n18500), .A2(n18906), .B1(n2465), .B2(n18908), .ZN(
        n3884) );
  OAI22_X1 U2866 ( .A1(n18497), .A2(n18905), .B1(n2456), .B2(n18908), .ZN(
        n3868) );
  OAI22_X1 U2867 ( .A1(n18494), .A2(n18906), .B1(n2447), .B2(n18908), .ZN(
        n3852) );
  OAI22_X1 U2868 ( .A1(n18491), .A2(n18905), .B1(n2438), .B2(n18908), .ZN(
        n3836) );
  OAI22_X1 U2869 ( .A1(n18442), .A2(n18740), .B1(n2281), .B2(n18743), .ZN(
        n2998) );
  OAI22_X1 U2870 ( .A1(n18439), .A2(n18741), .B1(n2272), .B2(n18743), .ZN(
        n2999) );
  OAI22_X1 U2871 ( .A1(n18436), .A2(n18740), .B1(n2263), .B2(n18743), .ZN(
        n3000) );
  OAI22_X1 U2872 ( .A1(n18433), .A2(n18741), .B1(n2254), .B2(n18743), .ZN(
        n3001) );
  OAI22_X1 U2873 ( .A1(n18430), .A2(n18740), .B1(n2245), .B2(n18742), .ZN(
        n3002) );
  OAI22_X1 U2874 ( .A1(n18427), .A2(n18741), .B1(n2236), .B2(n18742), .ZN(
        n3003) );
  OAI22_X1 U2875 ( .A1(n18424), .A2(n18740), .B1(n2227), .B2(n18742), .ZN(
        n3004) );
  OAI22_X1 U2876 ( .A1(n18421), .A2(n18741), .B1(n2218), .B2(n18742), .ZN(
        n3005) );
  OAI22_X1 U2877 ( .A1(n18440), .A2(n19015), .B1(n2286), .B2(n19018), .ZN(
        n9070) );
  OAI22_X1 U2878 ( .A1(n18437), .A2(n19016), .B1(n2277), .B2(n19018), .ZN(
        n9071) );
  OAI22_X1 U2879 ( .A1(n18434), .A2(n19015), .B1(n2268), .B2(n19018), .ZN(
        n9072) );
  OAI22_X1 U2880 ( .A1(n18431), .A2(n19016), .B1(n2259), .B2(n19018), .ZN(
        n9073) );
  OAI22_X1 U2881 ( .A1(n18428), .A2(n19015), .B1(n2250), .B2(n19017), .ZN(
        n9074) );
  OAI22_X1 U2882 ( .A1(n18425), .A2(n19016), .B1(n2241), .B2(n19017), .ZN(
        n9075) );
  OAI22_X1 U2883 ( .A1(n18422), .A2(n19015), .B1(n2232), .B2(n19017), .ZN(
        n9076) );
  OAI22_X1 U2884 ( .A1(n18419), .A2(n19016), .B1(n2223), .B2(n19017), .ZN(
        n9077) );
  NAND2_X1 U2885 ( .A1(n1753), .A2(n1754), .ZN(N1044) );
  NOR4_X1 U2886 ( .A1(n1763), .A2(n1764), .A3(n1765), .A4(n1766), .ZN(n1753)
         );
  NAND2_X1 U2887 ( .A1(n1735), .A2(n1736), .ZN(N1045) );
  NOR4_X1 U2888 ( .A1(n1745), .A2(n1746), .A3(n1747), .A4(n1748), .ZN(n1735)
         );
  NAND2_X1 U2889 ( .A1(n1717), .A2(n1718), .ZN(N1046) );
  NOR4_X1 U2890 ( .A1(n1727), .A2(n1728), .A3(n1729), .A4(n1730), .ZN(n1717)
         );
  NAND2_X1 U2891 ( .A1(n1699), .A2(n1700), .ZN(N1047) );
  NOR4_X1 U2892 ( .A1(n1709), .A2(n1710), .A3(n1711), .A4(n1712), .ZN(n1699)
         );
  NAND2_X1 U2893 ( .A1(n1681), .A2(n1682), .ZN(N1048) );
  NOR4_X1 U2894 ( .A1(n1691), .A2(n1692), .A3(n1693), .A4(n1694), .ZN(n1681)
         );
  NAND2_X1 U2895 ( .A1(n1663), .A2(n1664), .ZN(N1049) );
  NOR4_X1 U2896 ( .A1(n1673), .A2(n1674), .A3(n1675), .A4(n1676), .ZN(n1663)
         );
  NAND2_X1 U2897 ( .A1(n1645), .A2(n1646), .ZN(N1050) );
  NOR4_X1 U2898 ( .A1(n1655), .A2(n1656), .A3(n1657), .A4(n1658), .ZN(n1645)
         );
  NAND2_X1 U2899 ( .A1(n1595), .A2(n1596), .ZN(N1051) );
  NOR4_X1 U2900 ( .A1(n1621), .A2(n1622), .A3(n1623), .A4(n1624), .ZN(n1595)
         );
  AND3_X1 U2901 ( .A1(ADD_RD2[1]), .A2(n19920), .A3(ADD_RD2[2]), .ZN(n2194) );
  AND3_X1 U2902 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[0]), .A3(ADD_RD2[2]), .ZN(n2193) );
  INV_X1 U2903 ( .A(ADD_WR[0]), .ZN(n19126) );
  INV_X1 U2904 ( .A(ADD_WR[2]), .ZN(n19124) );
  INV_X1 U2905 ( .A(ADD_WR[1]), .ZN(n19125) );
  AND3_X1 U2906 ( .A1(n19920), .A2(n19921), .A3(ADD_RD2[2]), .ZN(n2196) );
  AND3_X1 U2907 ( .A1(ADD_RD2[0]), .A2(n19921), .A3(ADD_RD2[2]), .ZN(n2195) );
  INV_X1 U2908 ( .A(ADD_RD2[1]), .ZN(n19921) );
  INV_X1 U2909 ( .A(ADD_RD2[0]), .ZN(n19920) );
  NAND2_X1 U2910 ( .A1(n1259), .A2(n1260), .ZN(N707) );
  NOR4_X1 U2911 ( .A1(n1261), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1260)
         );
  NOR4_X1 U2912 ( .A1(n1269), .A2(n1270), .A3(n1271), .A4(n1272), .ZN(n1259)
         );
  OAI221_X1 U2913 ( .B1(n19757), .B2(n18669), .C1(n17973), .C2(n18666), .A(
        n1268), .ZN(n1261) );
  NAND2_X1 U2914 ( .A1(n1331), .A2(n1332), .ZN(N703) );
  NOR4_X1 U2915 ( .A1(n1333), .A2(n1334), .A3(n1335), .A4(n1336), .ZN(n1332)
         );
  NOR4_X1 U2916 ( .A1(n1341), .A2(n1342), .A3(n1343), .A4(n1344), .ZN(n1331)
         );
  OAI221_X1 U2917 ( .B1(n19761), .B2(n18669), .C1(n17969), .C2(n18666), .A(
        n1340), .ZN(n1333) );
  NAND2_X1 U2918 ( .A1(n1205), .A2(n1206), .ZN(N710) );
  NOR4_X1 U2919 ( .A1(n1207), .A2(n1208), .A3(n1209), .A4(n1210), .ZN(n1206)
         );
  NOR4_X1 U2920 ( .A1(n1215), .A2(n1216), .A3(n1217), .A4(n1218), .ZN(n1205)
         );
  OAI221_X1 U2921 ( .B1(n19754), .B2(n18669), .C1(n17976), .C2(n18666), .A(
        n1214), .ZN(n1207) );
  NAND2_X1 U2922 ( .A1(n1241), .A2(n1242), .ZN(N708) );
  NOR4_X1 U2923 ( .A1(n1243), .A2(n1244), .A3(n1245), .A4(n1246), .ZN(n1242)
         );
  NOR4_X1 U2924 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1241)
         );
  OAI221_X1 U2925 ( .B1(n19756), .B2(n18669), .C1(n17974), .C2(n18666), .A(
        n1250), .ZN(n1243) );
  NAND2_X1 U2926 ( .A1(n1313), .A2(n1314), .ZN(N704) );
  NOR4_X1 U2927 ( .A1(n1315), .A2(n1316), .A3(n1317), .A4(n1318), .ZN(n1314)
         );
  NOR4_X1 U2928 ( .A1(n1323), .A2(n1324), .A3(n1325), .A4(n1326), .ZN(n1313)
         );
  OAI221_X1 U2929 ( .B1(n19760), .B2(n18669), .C1(n17970), .C2(n18666), .A(
        n1322), .ZN(n1315) );
  NAND2_X1 U2930 ( .A1(n1187), .A2(n1188), .ZN(N711) );
  NOR4_X1 U2931 ( .A1(n1189), .A2(n1190), .A3(n1191), .A4(n1192), .ZN(n1188)
         );
  NOR4_X1 U2932 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1187)
         );
  OAI221_X1 U2933 ( .B1(n19753), .B2(n18669), .C1(n17977), .C2(n18666), .A(
        n1196), .ZN(n1189) );
  NAND2_X1 U2934 ( .A1(n1385), .A2(n1386), .ZN(N700) );
  NOR4_X1 U2935 ( .A1(n1387), .A2(n1388), .A3(n1389), .A4(n1390), .ZN(n1386)
         );
  NOR4_X1 U2936 ( .A1(n1395), .A2(n1396), .A3(n1397), .A4(n1398), .ZN(n1385)
         );
  OAI221_X1 U2937 ( .B1(n19764), .B2(n18668), .C1(n17966), .C2(n18665), .A(
        n1394), .ZN(n1387) );
  INV_X1 U2938 ( .A(ADD_RD1[0]), .ZN(n19914) );
  NAND2_X1 U2939 ( .A1(n1223), .A2(n1224), .ZN(N709) );
  NOR4_X1 U2940 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1224)
         );
  NOR4_X1 U2941 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .ZN(n1223)
         );
  OAI221_X1 U2942 ( .B1(n19755), .B2(n18669), .C1(n17975), .C2(n18666), .A(
        n1232), .ZN(n1225) );
  NAND2_X1 U2943 ( .A1(n1295), .A2(n1296), .ZN(N705) );
  NOR4_X1 U2944 ( .A1(n1297), .A2(n1298), .A3(n1299), .A4(n1300), .ZN(n1296)
         );
  NOR4_X1 U2945 ( .A1(n1305), .A2(n1306), .A3(n1307), .A4(n1308), .ZN(n1295)
         );
  OAI221_X1 U2946 ( .B1(n19759), .B2(n18669), .C1(n17971), .C2(n18666), .A(
        n1304), .ZN(n1297) );
  NAND2_X1 U2947 ( .A1(n1169), .A2(n1170), .ZN(N712) );
  NOR4_X1 U2948 ( .A1(n1171), .A2(n1172), .A3(n1173), .A4(n1174), .ZN(n1170)
         );
  NOR4_X1 U2949 ( .A1(n1179), .A2(n1180), .A3(n1181), .A4(n1182), .ZN(n1169)
         );
  OAI221_X1 U2950 ( .B1(n19752), .B2(n18669), .C1(n17978), .C2(n18666), .A(
        n1178), .ZN(n1171) );
  NAND2_X1 U2951 ( .A1(n1367), .A2(n1368), .ZN(N701) );
  NOR4_X1 U2952 ( .A1(n1369), .A2(n1370), .A3(n1371), .A4(n1372), .ZN(n1368)
         );
  NOR4_X1 U2953 ( .A1(n1377), .A2(n1378), .A3(n1379), .A4(n1380), .ZN(n1367)
         );
  OAI221_X1 U2954 ( .B1(n19763), .B2(n18668), .C1(n17967), .C2(n18665), .A(
        n1376), .ZN(n1369) );
  NAND2_X1 U2955 ( .A1(n1277), .A2(n1278), .ZN(N706) );
  NOR4_X1 U2956 ( .A1(n1279), .A2(n1280), .A3(n1281), .A4(n1282), .ZN(n1278)
         );
  NOR4_X1 U2957 ( .A1(n1287), .A2(n1288), .A3(n1289), .A4(n1290), .ZN(n1277)
         );
  OAI221_X1 U2958 ( .B1(n19758), .B2(n18669), .C1(n17972), .C2(n18666), .A(
        n1286), .ZN(n1279) );
  NAND2_X1 U2959 ( .A1(n1151), .A2(n1152), .ZN(N713) );
  NOR4_X1 U2960 ( .A1(n1153), .A2(n1154), .A3(n1155), .A4(n1156), .ZN(n1152)
         );
  NOR4_X1 U2961 ( .A1(n1161), .A2(n1162), .A3(n1163), .A4(n1164), .ZN(n1151)
         );
  OAI221_X1 U2962 ( .B1(n19751), .B2(n18669), .C1(n17979), .C2(n18666), .A(
        n1160), .ZN(n1153) );
  NAND2_X1 U2963 ( .A1(n1349), .A2(n1350), .ZN(N702) );
  NOR4_X1 U2964 ( .A1(n1351), .A2(n1352), .A3(n1353), .A4(n1354), .ZN(n1350)
         );
  NOR4_X1 U2965 ( .A1(n1359), .A2(n1360), .A3(n1361), .A4(n1362), .ZN(n1349)
         );
  OAI221_X1 U2966 ( .B1(n19762), .B2(n18669), .C1(n17968), .C2(n18666), .A(
        n1358), .ZN(n1351) );
  INV_X1 U2967 ( .A(ADD_RD1[1]), .ZN(n19917) );
  AND3_X1 U2968 ( .A1(ENABLE), .A2(n19057), .A3(WR), .ZN(n970) );
  NAND2_X1 U2969 ( .A1(n2185), .A2(n2186), .ZN(N1020) );
  NOR4_X1 U2970 ( .A1(n2187), .A2(n2188), .A3(n2189), .A4(n2190), .ZN(n2186)
         );
  NAND2_X1 U2971 ( .A1(n2167), .A2(n2168), .ZN(N1021) );
  NOR4_X1 U2972 ( .A1(n2169), .A2(n2170), .A3(n2171), .A4(n2172), .ZN(n2168)
         );
  NAND2_X1 U2973 ( .A1(n2149), .A2(n2150), .ZN(N1022) );
  NOR4_X1 U2974 ( .A1(n2151), .A2(n2152), .A3(n2153), .A4(n2154), .ZN(n2150)
         );
  NAND2_X1 U2975 ( .A1(n2131), .A2(n2132), .ZN(N1023) );
  NOR4_X1 U2976 ( .A1(n2133), .A2(n2134), .A3(n2135), .A4(n2136), .ZN(n2132)
         );
  NAND2_X1 U2977 ( .A1(n2113), .A2(n2114), .ZN(N1024) );
  NOR4_X1 U2978 ( .A1(n2115), .A2(n2116), .A3(n2117), .A4(n2118), .ZN(n2114)
         );
  NAND2_X1 U2979 ( .A1(n2095), .A2(n2096), .ZN(N1025) );
  NOR4_X1 U2980 ( .A1(n2097), .A2(n2098), .A3(n2099), .A4(n2100), .ZN(n2096)
         );
  NAND2_X1 U2981 ( .A1(n2077), .A2(n2078), .ZN(N1026) );
  NOR4_X1 U2982 ( .A1(n2079), .A2(n2080), .A3(n2081), .A4(n2082), .ZN(n2078)
         );
  INV_X1 U2983 ( .A(ADD_RD2[4]), .ZN(n19918) );
  INV_X1 U2984 ( .A(ADD_RD2[3]), .ZN(n19919) );
  INV_X1 U2985 ( .A(ADD_RD1[4]), .ZN(n19915) );
  INV_X1 U2986 ( .A(ADD_RD1[3]), .ZN(n19916) );
  NAND2_X1 U2987 ( .A1(n2059), .A2(n2060), .ZN(N1027) );
  NOR4_X1 U2988 ( .A1(n2061), .A2(n2062), .A3(n2063), .A4(n2064), .ZN(n2060)
         );
  NAND2_X1 U2989 ( .A1(n2041), .A2(n2042), .ZN(N1028) );
  NOR4_X1 U2990 ( .A1(n2051), .A2(n2052), .A3(n2053), .A4(n2054), .ZN(n2041)
         );
  NAND2_X1 U2991 ( .A1(n2023), .A2(n2024), .ZN(N1029) );
  NOR4_X1 U2992 ( .A1(n2033), .A2(n2034), .A3(n2035), .A4(n2036), .ZN(n2023)
         );
  NAND2_X1 U2993 ( .A1(n2005), .A2(n2006), .ZN(N1030) );
  NOR4_X1 U2994 ( .A1(n2015), .A2(n2016), .A3(n2017), .A4(n2018), .ZN(n2005)
         );
  NAND2_X1 U2995 ( .A1(n1987), .A2(n1988), .ZN(N1031) );
  NOR4_X1 U2996 ( .A1(n1997), .A2(n1998), .A3(n1999), .A4(n2000), .ZN(n1987)
         );
  NAND2_X1 U2997 ( .A1(n1969), .A2(n1970), .ZN(N1032) );
  NOR4_X1 U2998 ( .A1(n1979), .A2(n1980), .A3(n1981), .A4(n1982), .ZN(n1969)
         );
  NAND2_X1 U2999 ( .A1(n1951), .A2(n1952), .ZN(N1033) );
  NOR4_X1 U3000 ( .A1(n1961), .A2(n1962), .A3(n1963), .A4(n1964), .ZN(n1951)
         );
  NAND2_X1 U3001 ( .A1(n1933), .A2(n1934), .ZN(N1034) );
  NOR4_X1 U3002 ( .A1(n1943), .A2(n1944), .A3(n1945), .A4(n1946), .ZN(n1933)
         );
  NAND2_X1 U3003 ( .A1(n1915), .A2(n1916), .ZN(N1035) );
  NOR4_X1 U3004 ( .A1(n1925), .A2(n1926), .A3(n1927), .A4(n1928), .ZN(n1915)
         );
  NAND2_X1 U3005 ( .A1(n1897), .A2(n1898), .ZN(N1036) );
  NOR4_X1 U3006 ( .A1(n1907), .A2(n1908), .A3(n1909), .A4(n1910), .ZN(n1897)
         );
  NAND2_X1 U3007 ( .A1(n1879), .A2(n1880), .ZN(N1037) );
  NOR4_X1 U3008 ( .A1(n1889), .A2(n1890), .A3(n1891), .A4(n1892), .ZN(n1879)
         );
  NAND2_X1 U3009 ( .A1(n1861), .A2(n1862), .ZN(N1038) );
  NOR4_X1 U3010 ( .A1(n1871), .A2(n1872), .A3(n1873), .A4(n1874), .ZN(n1861)
         );
  NAND2_X1 U3011 ( .A1(n1843), .A2(n1844), .ZN(N1039) );
  NOR4_X1 U3012 ( .A1(n1853), .A2(n1854), .A3(n1855), .A4(n1856), .ZN(n1843)
         );
  NAND2_X1 U3013 ( .A1(n1825), .A2(n1826), .ZN(N1040) );
  NOR4_X1 U3014 ( .A1(n1835), .A2(n1836), .A3(n1837), .A4(n1838), .ZN(n1825)
         );
  NAND2_X1 U3015 ( .A1(n1807), .A2(n1808), .ZN(N1041) );
  NOR4_X1 U3016 ( .A1(n1817), .A2(n1818), .A3(n1819), .A4(n1820), .ZN(n1807)
         );
  NAND2_X1 U3017 ( .A1(n1789), .A2(n1790), .ZN(N1042) );
  NOR4_X1 U3018 ( .A1(n1799), .A2(n1800), .A3(n1801), .A4(n1802), .ZN(n1789)
         );
  NAND2_X1 U3019 ( .A1(n1771), .A2(n1772), .ZN(N1043) );
  NOR4_X1 U3020 ( .A1(n1781), .A2(n1782), .A3(n1783), .A4(n1784), .ZN(n1771)
         );
  INV_X1 U3021 ( .A(ADD_WR[4]), .ZN(n19122) );
  INV_X1 U3022 ( .A(ADD_WR[3]), .ZN(n19123) );
  INV_X1 U3023 ( .A(n903), .ZN(n19121) );
  AOI22_X1 U3024 ( .A1(DATAIN[0]), .A2(n19027), .B1(n19028), .B2(n17687), .ZN(
        n903) );
  INV_X1 U3025 ( .A(n905), .ZN(n19119) );
  AOI22_X1 U3026 ( .A1(DATAIN[1]), .A2(n19026), .B1(n19028), .B2(n17688), .ZN(
        n905) );
  INV_X1 U3027 ( .A(n906), .ZN(n19117) );
  AOI22_X1 U3028 ( .A1(DATAIN[2]), .A2(n19027), .B1(n19028), .B2(n17689), .ZN(
        n906) );
  INV_X1 U3029 ( .A(n907), .ZN(n19115) );
  AOI22_X1 U3030 ( .A1(DATAIN[3]), .A2(n19026), .B1(n19028), .B2(n17690), .ZN(
        n907) );
  INV_X1 U3031 ( .A(n908), .ZN(n19113) );
  AOI22_X1 U3032 ( .A1(DATAIN[4]), .A2(n19027), .B1(n19028), .B2(n17691), .ZN(
        n908) );
  INV_X1 U3033 ( .A(n909), .ZN(n19111) );
  AOI22_X1 U3034 ( .A1(DATAIN[5]), .A2(n19026), .B1(n19029), .B2(n17692), .ZN(
        n909) );
  INV_X1 U3035 ( .A(n910), .ZN(n19109) );
  AOI22_X1 U3036 ( .A1(DATAIN[6]), .A2(n19027), .B1(n19029), .B2(n17693), .ZN(
        n910) );
  INV_X1 U3037 ( .A(n911), .ZN(n19107) );
  AOI22_X1 U3038 ( .A1(DATAIN[7]), .A2(n19026), .B1(n19029), .B2(n17694), .ZN(
        n911) );
  INV_X1 U3039 ( .A(n912), .ZN(n19105) );
  AOI22_X1 U3040 ( .A1(DATAIN[8]), .A2(n19027), .B1(n19029), .B2(n17599), .ZN(
        n912) );
  INV_X1 U3041 ( .A(n913), .ZN(n19103) );
  AOI22_X1 U3042 ( .A1(DATAIN[9]), .A2(n19027), .B1(n19029), .B2(n17600), .ZN(
        n913) );
  INV_X1 U3043 ( .A(n914), .ZN(n19101) );
  AOI22_X1 U3044 ( .A1(DATAIN[10]), .A2(n19027), .B1(n19030), .B2(n17601), 
        .ZN(n914) );
  INV_X1 U3045 ( .A(n915), .ZN(n19099) );
  AOI22_X1 U3046 ( .A1(DATAIN[11]), .A2(n19027), .B1(n19030), .B2(n17602), 
        .ZN(n915) );
  INV_X1 U3047 ( .A(n916), .ZN(n19097) );
  AOI22_X1 U3048 ( .A1(DATAIN[12]), .A2(n19027), .B1(n19030), .B2(n17603), 
        .ZN(n916) );
  INV_X1 U3049 ( .A(n917), .ZN(n19095) );
  AOI22_X1 U3050 ( .A1(DATAIN[13]), .A2(n19027), .B1(n19030), .B2(n17604), 
        .ZN(n917) );
  INV_X1 U3051 ( .A(n918), .ZN(n19093) );
  AOI22_X1 U3052 ( .A1(DATAIN[14]), .A2(n19027), .B1(n19030), .B2(n17605), 
        .ZN(n918) );
  INV_X1 U3053 ( .A(n919), .ZN(n19091) );
  AOI22_X1 U3054 ( .A1(DATAIN[15]), .A2(n19027), .B1(n19031), .B2(n17606), 
        .ZN(n919) );
  INV_X1 U3055 ( .A(n920), .ZN(n19089) );
  AOI22_X1 U3056 ( .A1(DATAIN[16]), .A2(n19027), .B1(n19031), .B2(n17607), 
        .ZN(n920) );
  INV_X1 U3057 ( .A(n921), .ZN(n19087) );
  AOI22_X1 U3058 ( .A1(DATAIN[17]), .A2(n19027), .B1(n19031), .B2(n17608), 
        .ZN(n921) );
  INV_X1 U3059 ( .A(n922), .ZN(n19085) );
  AOI22_X1 U3060 ( .A1(DATAIN[18]), .A2(n19027), .B1(n19031), .B2(n17609), 
        .ZN(n922) );
  INV_X1 U3061 ( .A(n923), .ZN(n19083) );
  AOI22_X1 U3062 ( .A1(DATAIN[19]), .A2(n19027), .B1(n19031), .B2(n17610), 
        .ZN(n923) );
  INV_X1 U3063 ( .A(n924), .ZN(n19081) );
  AOI22_X1 U3064 ( .A1(DATAIN[20]), .A2(n19026), .B1(n19032), .B2(n17611), 
        .ZN(n924) );
  INV_X1 U3065 ( .A(n925), .ZN(n19079) );
  AOI22_X1 U3066 ( .A1(DATAIN[21]), .A2(n19026), .B1(n19032), .B2(n17612), 
        .ZN(n925) );
  INV_X1 U3067 ( .A(n926), .ZN(n19077) );
  AOI22_X1 U3068 ( .A1(DATAIN[22]), .A2(n19026), .B1(n19032), .B2(n17613), 
        .ZN(n926) );
  INV_X1 U3069 ( .A(n927), .ZN(n19075) );
  AOI22_X1 U3070 ( .A1(DATAIN[23]), .A2(n19026), .B1(n19032), .B2(n17614), 
        .ZN(n927) );
  INV_X1 U3071 ( .A(n928), .ZN(n19073) );
  AOI22_X1 U3072 ( .A1(DATAIN[24]), .A2(n19026), .B1(n19032), .B2(n17615), 
        .ZN(n928) );
  INV_X1 U3073 ( .A(n929), .ZN(n19071) );
  AOI22_X1 U3074 ( .A1(DATAIN[25]), .A2(n19026), .B1(n19033), .B2(n17616), 
        .ZN(n929) );
  INV_X1 U3075 ( .A(n930), .ZN(n19069) );
  AOI22_X1 U3076 ( .A1(DATAIN[26]), .A2(n19026), .B1(n19033), .B2(n17617), 
        .ZN(n930) );
  INV_X1 U3077 ( .A(n931), .ZN(n19067) );
  AOI22_X1 U3078 ( .A1(DATAIN[27]), .A2(n19026), .B1(n19033), .B2(n17618), 
        .ZN(n931) );
  INV_X1 U3079 ( .A(n932), .ZN(n19065) );
  AOI22_X1 U3080 ( .A1(DATAIN[28]), .A2(n19026), .B1(n19033), .B2(n17619), 
        .ZN(n932) );
  INV_X1 U3081 ( .A(n933), .ZN(n19063) );
  AOI22_X1 U3082 ( .A1(DATAIN[29]), .A2(n19026), .B1(n19033), .B2(n17620), 
        .ZN(n933) );
  INV_X1 U3083 ( .A(n934), .ZN(n19061) );
  AOI22_X1 U3084 ( .A1(DATAIN[30]), .A2(n19026), .B1(n19034), .B2(n17621), 
        .ZN(n934) );
  INV_X1 U3085 ( .A(n935), .ZN(n19059) );
  AOI22_X1 U3086 ( .A1(DATAIN[31]), .A2(n19026), .B1(n19034), .B2(n17622), 
        .ZN(n935) );
  NOR3_X1 U3087 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n19914), .ZN(n1577) );
  NOR3_X1 U3088 ( .A1(n19914), .A2(ADD_RD1[2]), .A3(n19917), .ZN(n1579) );
  NOR3_X1 U3089 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(ADD_RD1[0]), .ZN(n1576) );
  OAI221_X1 U3090 ( .B1(n17877), .B2(n18656), .C1(n18177), .C2(n18653), .A(
        n1471), .ZN(n1470) );
  NOR3_X1 U3091 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[2]), .A3(n19917), .ZN(n1572) );
endmodule


module DecodeUnit_DW01_add_0 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [9:1] carry;

  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XOR2_X1 U3 ( .A(A[6]), .B(B[6]), .Z(n3) );
  XOR2_X1 U4 ( .A(n3), .B(carry[6]), .Z(SUM[6]) );
  NAND3_X1 U8 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[7]) );
  XOR2_X1 U9 ( .A(A[7]), .B(B[7]), .Z(n7) );
  XOR2_X1 U10 ( .A(n7), .B(carry[7]), .Z(SUM[7]) );
  NAND3_X1 U14 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[8]) );
  XOR2_X1 U15 ( .A(B[1]), .B(A[1]), .Z(n11) );
  XOR2_X1 U16 ( .A(n2), .B(n11), .Z(SUM[1]) );
  NAND3_X1 U20 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[2]) );
  XOR2_X1 U21 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR2_X1 U22 ( .A(carry[2]), .B(n15), .Z(SUM[2]) );
  NAND3_X1 U26 ( .A1(n16), .A2(n17), .A3(n18), .ZN(carry[3]) );
  XOR2_X1 U27 ( .A(B[9]), .B(A[9]), .Z(n19) );
  XOR2_X1 U28 ( .A(carry[9]), .B(n19), .Z(SUM[9]) );
  NAND2_X1 U2 ( .A1(A[6]), .A2(B[6]), .ZN(n4) );
  NAND2_X1 U5 ( .A1(A[6]), .A2(carry[6]), .ZN(n5) );
  NAND2_X1 U6 ( .A1(B[6]), .A2(carry[6]), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n2), .A2(B[1]), .ZN(n12) );
  NAND2_X1 U11 ( .A1(n2), .A2(A[1]), .ZN(n13) );
  NAND2_X1 U12 ( .A1(B[1]), .A2(A[1]), .ZN(n14) );
  NAND2_X1 U13 ( .A1(B[2]), .A2(A[2]), .ZN(n18) );
  NAND2_X1 U17 ( .A1(carry[2]), .A2(B[2]), .ZN(n16) );
  AND2_X1 U18 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
  NAND2_X1 U19 ( .A1(A[7]), .A2(B[7]), .ZN(n8) );
  NAND2_X1 U23 ( .A1(A[7]), .A2(carry[7]), .ZN(n9) );
  NAND2_X1 U24 ( .A1(B[7]), .A2(carry[7]), .ZN(n10) );
  NAND2_X1 U25 ( .A1(carry[2]), .A2(A[2]), .ZN(n17) );
endmodule


module DecodeUnit ( clock, reset, JMP, RegDestination, en2, SignSelect, 
        BranchCondSel, BRANCHenable, RD1, RD2, WR, Instruction, ADD_WR, DATAIN, 
        NPCfromIF, OUT1, OUT2, OUTNPC, OUTIMM, NPCtoEX, AddressWtoEX, 
        BRANCHtoFetch );
  input [31:0] Instruction;
  input [4:0] ADD_WR;
  input [31:0] DATAIN;
  input [31:0] NPCfromIF;
  output [31:0] OUT1;
  output [31:0] OUT2;
  output [31:0] OUTNPC;
  output [31:0] OUTIMM;
  output [31:0] NPCtoEX;
  output [31:0] AddressWtoEX;
  input clock, reset, JMP, RegDestination, en2, SignSelect, BranchCondSel,
         BRANCHenable, RD1, RD2, WR;
  output BRANCHtoFetch;
  wire   BranchTaken, n4;
  wire   [31:0] AddressW;
  wire   [31:0] MuxtoIMM;
  wire   [31:0] RFOUT1;
  wire   [31:0] RFOUT2;
  assign OUTNPC[10] = 1'b0;
  assign OUTNPC[11] = 1'b0;
  assign OUTNPC[12] = 1'b0;
  assign OUTNPC[13] = 1'b0;
  assign OUTNPC[14] = 1'b0;
  assign OUTNPC[15] = 1'b0;
  assign OUTNPC[16] = 1'b0;
  assign OUTNPC[17] = 1'b0;
  assign OUTNPC[18] = 1'b0;
  assign OUTNPC[19] = 1'b0;
  assign OUTNPC[20] = 1'b0;
  assign OUTNPC[21] = 1'b0;
  assign OUTNPC[22] = 1'b0;
  assign OUTNPC[23] = 1'b0;
  assign OUTNPC[24] = 1'b0;
  assign OUTNPC[25] = 1'b0;
  assign OUTNPC[26] = 1'b0;
  assign OUTNPC[27] = 1'b0;
  assign OUTNPC[28] = 1'b0;
  assign OUTNPC[29] = 1'b0;
  assign OUTNPC[30] = 1'b0;
  assign OUTNPC[31] = 1'b0;

  Mux41 ADDRESS_MUX ( .a({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Instruction[20:16]}), .b({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, Instruction[15:11]}), .c({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1}), .d({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .sel({JMP, RegDestination}), .y(AddressW) );
  Mux21_5 MUX ( .a({Instruction[15], Instruction[15], Instruction[15], 
        Instruction[15], Instruction[15], Instruction[15], Instruction[15], 
        Instruction[15], Instruction[15], Instruction[15], Instruction[15], 
        Instruction[15], Instruction[15], Instruction[15], Instruction[15], 
        Instruction[15], Instruction[15:0]}), .b({Instruction[25], 
        Instruction[25], Instruction[25], Instruction[25], Instruction[25], 
        Instruction[25], Instruction[25:0]}), .sel(SignSelect), .y(MuxtoIMM)
         );
  BranchUnit BRANCH ( .a(RFOUT1), .sel(BranchCondSel), .y(BranchTaken) );
  reg_11 IMM_REG ( .clock(clock), .reset(reset), .load(en2), .i(MuxtoIMM), .o(
        OUTIMM) );
  reg_10 OUT1_REG ( .clock(clock), .reset(reset), .load(en2), .i(RFOUT1), .o(
        OUT1) );
  reg_9 OUT2_REG ( .clock(clock), .reset(reset), .load(en2), .i(RFOUT2), .o(
        OUT2) );
  reg_8 NXPC_REG ( .clock(clock), .reset(reset), .load(en2), .i(NPCfromIF), 
        .o(NPCtoEX) );
  reg_7 ADD_WR_REG ( .clock(clock), .reset(reset), .load(en2), .i(AddressW), 
        .o(AddressWtoEX) );
  register_file RF ( .CLK(clock), .RESET(reset), .ENABLE(1'b1), .RD1(RD1), 
        .RD2(RD2), .WR(WR), .ADD_WR(ADD_WR), .ADD_RD1(Instruction[25:21]), 
        .ADD_RD2(Instruction[20:16]), .DATAIN(DATAIN), .OUT1(RFOUT1), .OUT2(
        RFOUT2) );
  DecodeUnit_DW01_add_0 add_142 ( .A(NPCfromIF[9:0]), .B(MuxtoIMM[11:2]), .CI(
        1'b0), .SUM(OUTNPC[9:0]) );
  INV_X1 U3 ( .A(n4), .ZN(BRANCHtoFetch) );
  AOI21_X1 U5 ( .B1(BranchTaken), .B2(BRANCHenable), .A(JMP), .ZN(n4) );
endmodule


module Mux21_4 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397;

  INV_X1 U1 ( .A(n396), .ZN(n387) );
  BUF_X1 U2 ( .A(n397), .Z(n392) );
  BUF_X1 U3 ( .A(n397), .Z(n391) );
  BUF_X1 U4 ( .A(n397), .Z(n388) );
  BUF_X1 U5 ( .A(n397), .Z(n390) );
  BUF_X1 U6 ( .A(n397), .Z(n393) );
  BUF_X1 U7 ( .A(n388), .Z(n394) );
  BUF_X1 U8 ( .A(n389), .Z(n395) );
  BUF_X1 U9 ( .A(n397), .Z(n389) );
  BUF_X1 U10 ( .A(n392), .Z(n396) );
  INV_X1 U11 ( .A(n386), .ZN(n397) );
  INV_X1 U12 ( .A(n41), .ZN(y[31]) );
  AOI22_X1 U13 ( .A1(a[31]), .A2(sel), .B1(b[31]), .B2(n389), .ZN(n41) );
  INV_X1 U14 ( .A(n35), .ZN(y[8]) );
  AOI22_X1 U15 ( .A1(a[8]), .A2(n386), .B1(b[8]), .B2(n388), .ZN(n35) );
  INV_X1 U16 ( .A(n61), .ZN(y[13]) );
  AOI22_X1 U17 ( .A1(a[13]), .A2(n387), .B1(b[13]), .B2(n394), .ZN(n61) );
  INV_X1 U18 ( .A(n36), .ZN(y[7]) );
  AOI22_X1 U19 ( .A1(a[7]), .A2(sel), .B1(b[7]), .B2(n388), .ZN(n36) );
  INV_X1 U20 ( .A(n34), .ZN(y[9]) );
  AOI22_X1 U21 ( .A1(n386), .A2(a[9]), .B1(b[9]), .B2(n388), .ZN(n34) );
  INV_X1 U22 ( .A(n64), .ZN(y[10]) );
  AOI22_X1 U23 ( .A1(a[10]), .A2(n387), .B1(b[10]), .B2(n395), .ZN(n64) );
  INV_X1 U24 ( .A(n62), .ZN(y[12]) );
  AOI22_X1 U25 ( .A1(a[12]), .A2(n387), .B1(b[12]), .B2(n395), .ZN(n62) );
  INV_X1 U26 ( .A(n63), .ZN(y[11]) );
  AOI22_X1 U27 ( .A1(a[11]), .A2(n387), .B1(b[11]), .B2(n395), .ZN(n63) );
  INV_X1 U28 ( .A(n42), .ZN(y[30]) );
  AOI22_X1 U29 ( .A1(a[30]), .A2(sel), .B1(b[30]), .B2(n390), .ZN(n42) );
  INV_X1 U30 ( .A(n52), .ZN(y[21]) );
  AOI22_X1 U31 ( .A1(a[21]), .A2(n386), .B1(b[21]), .B2(n392), .ZN(n52) );
  INV_X1 U32 ( .A(n53), .ZN(y[20]) );
  AOI22_X1 U33 ( .A1(a[20]), .A2(sel), .B1(b[20]), .B2(n392), .ZN(n53) );
  INV_X1 U34 ( .A(n51), .ZN(y[22]) );
  AOI22_X1 U35 ( .A1(a[22]), .A2(n386), .B1(b[22]), .B2(n392), .ZN(n51) );
  INV_X1 U36 ( .A(n44), .ZN(y[29]) );
  AOI22_X1 U37 ( .A1(a[29]), .A2(sel), .B1(b[29]), .B2(n390), .ZN(n44) );
  INV_X1 U38 ( .A(n57), .ZN(y[17]) );
  AOI22_X1 U39 ( .A1(a[17]), .A2(n387), .B1(b[17]), .B2(n393), .ZN(n57) );
  INV_X1 U40 ( .A(n50), .ZN(y[23]) );
  AOI22_X1 U41 ( .A1(a[23]), .A2(n386), .B1(b[23]), .B2(n392), .ZN(n50) );
  INV_X1 U42 ( .A(n55), .ZN(y[19]) );
  AOI22_X1 U43 ( .A1(a[19]), .A2(n387), .B1(b[19]), .B2(n393), .ZN(n55) );
  INV_X1 U44 ( .A(n56), .ZN(y[18]) );
  AOI22_X1 U45 ( .A1(a[18]), .A2(n387), .B1(b[18]), .B2(n393), .ZN(n56) );
  INV_X1 U46 ( .A(n58), .ZN(y[16]) );
  AOI22_X1 U47 ( .A1(a[16]), .A2(n387), .B1(b[16]), .B2(n394), .ZN(n58) );
  INV_X1 U48 ( .A(n45), .ZN(y[28]) );
  AOI22_X1 U49 ( .A1(a[28]), .A2(sel), .B1(b[28]), .B2(n390), .ZN(n45) );
  INV_X1 U50 ( .A(n59), .ZN(y[15]) );
  AOI22_X1 U51 ( .A1(a[15]), .A2(n387), .B1(b[15]), .B2(n394), .ZN(n59) );
  INV_X1 U52 ( .A(n60), .ZN(y[14]) );
  AOI22_X1 U53 ( .A1(a[14]), .A2(n387), .B1(b[14]), .B2(n394), .ZN(n60) );
  INV_X1 U54 ( .A(n48), .ZN(y[25]) );
  AOI22_X1 U55 ( .A1(a[25]), .A2(n386), .B1(b[25]), .B2(n391), .ZN(n48) );
  INV_X1 U56 ( .A(n49), .ZN(y[24]) );
  AOI22_X1 U57 ( .A1(a[24]), .A2(sel), .B1(b[24]), .B2(n391), .ZN(n49) );
  INV_X1 U58 ( .A(n65), .ZN(y[0]) );
  AOI22_X1 U59 ( .A1(a[0]), .A2(n387), .B1(b[0]), .B2(n395), .ZN(n65) );
  INV_X1 U60 ( .A(n46), .ZN(y[27]) );
  AOI22_X1 U61 ( .A1(a[27]), .A2(n386), .B1(b[27]), .B2(n391), .ZN(n46) );
  INV_X1 U62 ( .A(n47), .ZN(y[26]) );
  AOI22_X1 U63 ( .A1(a[26]), .A2(sel), .B1(b[26]), .B2(n391), .ZN(n47) );
  INV_X1 U64 ( .A(n37), .ZN(y[6]) );
  AOI22_X1 U65 ( .A1(a[6]), .A2(n386), .B1(b[6]), .B2(n388), .ZN(n37) );
  INV_X1 U66 ( .A(n54), .ZN(y[1]) );
  AOI22_X1 U67 ( .A1(a[1]), .A2(n387), .B1(b[1]), .B2(n393), .ZN(n54) );
  INV_X1 U68 ( .A(n38), .ZN(y[5]) );
  AOI22_X1 U69 ( .A1(a[5]), .A2(sel), .B1(b[5]), .B2(n389), .ZN(n38) );
  INV_X1 U70 ( .A(n43), .ZN(y[2]) );
  AOI22_X1 U71 ( .A1(a[2]), .A2(n386), .B1(b[2]), .B2(n390), .ZN(n43) );
  INV_X1 U72 ( .A(n40), .ZN(y[3]) );
  AOI22_X1 U73 ( .A1(a[3]), .A2(n386), .B1(b[3]), .B2(n389), .ZN(n40) );
  INV_X1 U74 ( .A(n39), .ZN(y[4]) );
  AOI22_X1 U75 ( .A1(a[4]), .A2(sel), .B1(b[4]), .B2(n389), .ZN(n39) );
  BUF_X1 U76 ( .A(sel), .Z(n386) );
endmodule


module Mux21_3 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463;

  INV_X1 U1 ( .A(n398), .ZN(n388) );
  INV_X1 U2 ( .A(n398), .ZN(n387) );
  BUF_X1 U3 ( .A(n399), .Z(n392) );
  BUF_X1 U4 ( .A(n399), .Z(n397) );
  BUF_X1 U5 ( .A(n398), .Z(n396) );
  BUF_X1 U6 ( .A(n399), .Z(n395) );
  BUF_X1 U7 ( .A(n399), .Z(n394) );
  BUF_X1 U8 ( .A(n399), .Z(n393) );
  BUF_X1 U9 ( .A(n398), .Z(n391) );
  BUF_X1 U10 ( .A(n397), .Z(n390) );
  BUF_X1 U11 ( .A(n399), .Z(n398) );
  INV_X1 U12 ( .A(n386), .ZN(n399) );
  INV_X1 U13 ( .A(n455), .ZN(y[30]) );
  AOI22_X1 U14 ( .A1(a[30]), .A2(n388), .B1(b[30]), .B2(n392), .ZN(n455) );
  INV_X1 U15 ( .A(n453), .ZN(y[29]) );
  AOI22_X1 U16 ( .A1(a[29]), .A2(n388), .B1(b[29]), .B2(n392), .ZN(n453) );
  INV_X1 U17 ( .A(n449), .ZN(y[25]) );
  AOI22_X1 U18 ( .A1(a[25]), .A2(n388), .B1(b[25]), .B2(n393), .ZN(n449) );
  INV_X1 U19 ( .A(n438), .ZN(y[15]) );
  AOI22_X1 U20 ( .A1(a[15]), .A2(n387), .B1(b[15]), .B2(n396), .ZN(n438) );
  INV_X1 U21 ( .A(n448), .ZN(y[24]) );
  AOI22_X1 U22 ( .A1(a[24]), .A2(n388), .B1(b[24]), .B2(n393), .ZN(n448) );
  INV_X1 U23 ( .A(n456), .ZN(y[31]) );
  AOI22_X1 U24 ( .A1(a[31]), .A2(n389), .B1(b[31]), .B2(n391), .ZN(n456) );
  INV_X1 U25 ( .A(n436), .ZN(y[13]) );
  AOI22_X1 U26 ( .A1(a[13]), .A2(n387), .B1(b[13]), .B2(n396), .ZN(n436) );
  INV_X1 U27 ( .A(n446), .ZN(y[22]) );
  AOI22_X1 U28 ( .A1(a[22]), .A2(n388), .B1(b[22]), .B2(n394), .ZN(n446) );
  INV_X1 U29 ( .A(n452), .ZN(y[28]) );
  AOI22_X1 U30 ( .A1(a[28]), .A2(n388), .B1(b[28]), .B2(n392), .ZN(n452) );
  INV_X1 U31 ( .A(n435), .ZN(y[12]) );
  AOI22_X1 U32 ( .A1(a[12]), .A2(n387), .B1(b[12]), .B2(n397), .ZN(n435) );
  INV_X1 U33 ( .A(n450), .ZN(y[26]) );
  AOI22_X1 U34 ( .A1(a[26]), .A2(n388), .B1(b[26]), .B2(n393), .ZN(n450) );
  INV_X1 U35 ( .A(n447), .ZN(y[23]) );
  AOI22_X1 U36 ( .A1(a[23]), .A2(n388), .B1(b[23]), .B2(n394), .ZN(n447) );
  INV_X1 U37 ( .A(n440), .ZN(y[17]) );
  AOI22_X1 U38 ( .A1(a[17]), .A2(n387), .B1(b[17]), .B2(n395), .ZN(n440) );
  INV_X1 U39 ( .A(n463), .ZN(y[9]) );
  AOI22_X1 U40 ( .A1(n389), .A2(a[9]), .B1(b[9]), .B2(n390), .ZN(n463) );
  INV_X1 U41 ( .A(n462), .ZN(y[8]) );
  AOI22_X1 U42 ( .A1(a[8]), .A2(n389), .B1(b[8]), .B2(n390), .ZN(n462) );
  INV_X1 U43 ( .A(n439), .ZN(y[16]) );
  AOI22_X1 U44 ( .A1(a[16]), .A2(n387), .B1(b[16]), .B2(n396), .ZN(n439) );
  INV_X1 U45 ( .A(n444), .ZN(y[20]) );
  AOI22_X1 U46 ( .A1(a[20]), .A2(n388), .B1(b[20]), .B2(n394), .ZN(n444) );
  INV_X1 U47 ( .A(n434), .ZN(y[11]) );
  AOI22_X1 U48 ( .A1(a[11]), .A2(n387), .B1(b[11]), .B2(n397), .ZN(n434) );
  INV_X1 U49 ( .A(n442), .ZN(y[19]) );
  AOI22_X1 U50 ( .A1(a[19]), .A2(n387), .B1(b[19]), .B2(n395), .ZN(n442) );
  INV_X1 U51 ( .A(n451), .ZN(y[27]) );
  AOI22_X1 U52 ( .A1(a[27]), .A2(n388), .B1(b[27]), .B2(n393), .ZN(n451) );
  INV_X1 U53 ( .A(n433), .ZN(y[10]) );
  AOI22_X1 U54 ( .A1(a[10]), .A2(n387), .B1(b[10]), .B2(n397), .ZN(n433) );
  INV_X1 U55 ( .A(n437), .ZN(y[14]) );
  AOI22_X1 U56 ( .A1(a[14]), .A2(n387), .B1(b[14]), .B2(n396), .ZN(n437) );
  INV_X1 U57 ( .A(n441), .ZN(y[18]) );
  AOI22_X1 U58 ( .A1(a[18]), .A2(n387), .B1(b[18]), .B2(n395), .ZN(n441) );
  INV_X1 U59 ( .A(n445), .ZN(y[21]) );
  AOI22_X1 U60 ( .A1(a[21]), .A2(n388), .B1(b[21]), .B2(n394), .ZN(n445) );
  INV_X1 U61 ( .A(n443), .ZN(y[1]) );
  AOI22_X1 U62 ( .A1(a[1]), .A2(n387), .B1(b[1]), .B2(n395), .ZN(n443) );
  INV_X1 U63 ( .A(n454), .ZN(y[2]) );
  AOI22_X1 U64 ( .A1(a[2]), .A2(n388), .B1(b[2]), .B2(n392), .ZN(n454) );
  INV_X1 U65 ( .A(n458), .ZN(y[4]) );
  AOI22_X1 U66 ( .A1(a[4]), .A2(n389), .B1(b[4]), .B2(n391), .ZN(n458) );
  INV_X1 U67 ( .A(n459), .ZN(y[5]) );
  AOI22_X1 U68 ( .A1(a[5]), .A2(n389), .B1(b[5]), .B2(n391), .ZN(n459) );
  INV_X1 U69 ( .A(n460), .ZN(y[6]) );
  AOI22_X1 U70 ( .A1(a[6]), .A2(n389), .B1(b[6]), .B2(n390), .ZN(n460) );
  INV_X1 U71 ( .A(n461), .ZN(y[7]) );
  AOI22_X1 U72 ( .A1(a[7]), .A2(n389), .B1(b[7]), .B2(n390), .ZN(n461) );
  INV_X1 U73 ( .A(n457), .ZN(y[3]) );
  AOI22_X1 U74 ( .A1(a[3]), .A2(n389), .B1(b[3]), .B2(n391), .ZN(n457) );
  INV_X1 U75 ( .A(n432), .ZN(y[0]) );
  AOI22_X1 U76 ( .A1(a[0]), .A2(n387), .B1(b[0]), .B2(n397), .ZN(n432) );
  BUF_X1 U77 ( .A(sel), .Z(n386) );
  INV_X1 U78 ( .A(n398), .ZN(n389) );
endmodule


module Mux21_2 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462;

  INV_X1 U1 ( .A(n455), .ZN(y[31]) );
  INV_X1 U2 ( .A(n397), .ZN(n387) );
  INV_X1 U3 ( .A(n397), .ZN(n388) );
  BUF_X1 U4 ( .A(n398), .Z(n395) );
  BUF_X1 U5 ( .A(n398), .Z(n393) );
  BUF_X1 U6 ( .A(n397), .Z(n392) );
  BUF_X1 U7 ( .A(n398), .Z(n391) );
  BUF_X1 U8 ( .A(n397), .Z(n389) );
  BUF_X1 U9 ( .A(n398), .Z(n396) );
  BUF_X1 U10 ( .A(n398), .Z(n390) );
  BUF_X1 U11 ( .A(n391), .Z(n394) );
  BUF_X1 U12 ( .A(n398), .Z(n397) );
  INV_X1 U13 ( .A(n386), .ZN(n398) );
  AOI22_X1 U14 ( .A1(a[31]), .A2(n386), .B1(b[31]), .B2(n390), .ZN(n455) );
  INV_X1 U15 ( .A(n461), .ZN(y[8]) );
  AOI22_X1 U16 ( .A1(a[8]), .A2(sel), .B1(b[8]), .B2(n389), .ZN(n461) );
  INV_X1 U17 ( .A(n435), .ZN(y[13]) );
  AOI22_X1 U18 ( .A1(a[13]), .A2(n387), .B1(b[13]), .B2(n395), .ZN(n435) );
  INV_X1 U19 ( .A(n460), .ZN(y[7]) );
  AOI22_X1 U20 ( .A1(a[7]), .A2(n386), .B1(b[7]), .B2(n389), .ZN(n460) );
  INV_X1 U21 ( .A(n462), .ZN(y[9]) );
  AOI22_X1 U22 ( .A1(sel), .A2(a[9]), .B1(b[9]), .B2(n389), .ZN(n462) );
  INV_X1 U23 ( .A(n432), .ZN(y[10]) );
  AOI22_X1 U24 ( .A1(a[10]), .A2(n387), .B1(b[10]), .B2(n396), .ZN(n432) );
  INV_X1 U25 ( .A(n434), .ZN(y[12]) );
  AOI22_X1 U26 ( .A1(a[12]), .A2(n387), .B1(b[12]), .B2(n396), .ZN(n434) );
  INV_X1 U27 ( .A(n433), .ZN(y[11]) );
  AOI22_X1 U28 ( .A1(a[11]), .A2(n387), .B1(b[11]), .B2(n396), .ZN(n433) );
  INV_X1 U29 ( .A(n454), .ZN(y[30]) );
  AOI22_X1 U30 ( .A1(a[30]), .A2(n388), .B1(b[30]), .B2(n391), .ZN(n454) );
  INV_X1 U31 ( .A(n444), .ZN(y[21]) );
  AOI22_X1 U32 ( .A1(a[21]), .A2(n388), .B1(b[21]), .B2(n393), .ZN(n444) );
  INV_X1 U33 ( .A(n443), .ZN(y[20]) );
  AOI22_X1 U34 ( .A1(a[20]), .A2(n388), .B1(b[20]), .B2(n393), .ZN(n443) );
  INV_X1 U35 ( .A(n445), .ZN(y[22]) );
  AOI22_X1 U36 ( .A1(a[22]), .A2(n388), .B1(b[22]), .B2(n393), .ZN(n445) );
  INV_X1 U37 ( .A(n452), .ZN(y[29]) );
  AOI22_X1 U38 ( .A1(a[29]), .A2(n388), .B1(b[29]), .B2(n391), .ZN(n452) );
  INV_X1 U39 ( .A(n439), .ZN(y[17]) );
  AOI22_X1 U40 ( .A1(a[17]), .A2(n387), .B1(b[17]), .B2(n394), .ZN(n439) );
  INV_X1 U41 ( .A(n446), .ZN(y[23]) );
  AOI22_X1 U42 ( .A1(a[23]), .A2(n388), .B1(b[23]), .B2(n393), .ZN(n446) );
  INV_X1 U43 ( .A(n441), .ZN(y[19]) );
  AOI22_X1 U44 ( .A1(a[19]), .A2(n387), .B1(b[19]), .B2(n394), .ZN(n441) );
  INV_X1 U45 ( .A(n440), .ZN(y[18]) );
  AOI22_X1 U46 ( .A1(a[18]), .A2(n387), .B1(b[18]), .B2(n394), .ZN(n440) );
  INV_X1 U47 ( .A(n438), .ZN(y[16]) );
  AOI22_X1 U48 ( .A1(a[16]), .A2(n387), .B1(b[16]), .B2(n395), .ZN(n438) );
  INV_X1 U49 ( .A(n451), .ZN(y[28]) );
  AOI22_X1 U50 ( .A1(a[28]), .A2(n388), .B1(b[28]), .B2(n391), .ZN(n451) );
  INV_X1 U51 ( .A(n437), .ZN(y[15]) );
  AOI22_X1 U52 ( .A1(a[15]), .A2(n387), .B1(b[15]), .B2(n395), .ZN(n437) );
  INV_X1 U53 ( .A(n436), .ZN(y[14]) );
  AOI22_X1 U54 ( .A1(a[14]), .A2(n387), .B1(b[14]), .B2(n395), .ZN(n436) );
  INV_X1 U55 ( .A(n448), .ZN(y[25]) );
  AOI22_X1 U56 ( .A1(a[25]), .A2(n388), .B1(b[25]), .B2(n392), .ZN(n448) );
  INV_X1 U57 ( .A(n447), .ZN(y[24]) );
  AOI22_X1 U58 ( .A1(a[24]), .A2(n388), .B1(b[24]), .B2(n392), .ZN(n447) );
  INV_X1 U59 ( .A(n431), .ZN(y[0]) );
  AOI22_X1 U60 ( .A1(a[0]), .A2(n387), .B1(b[0]), .B2(n396), .ZN(n431) );
  INV_X1 U61 ( .A(n450), .ZN(y[27]) );
  AOI22_X1 U62 ( .A1(a[27]), .A2(n388), .B1(b[27]), .B2(n392), .ZN(n450) );
  INV_X1 U63 ( .A(n449), .ZN(y[26]) );
  AOI22_X1 U64 ( .A1(a[26]), .A2(n388), .B1(b[26]), .B2(n392), .ZN(n449) );
  INV_X1 U65 ( .A(n459), .ZN(y[6]) );
  AOI22_X1 U66 ( .A1(a[6]), .A2(sel), .B1(b[6]), .B2(n389), .ZN(n459) );
  INV_X1 U67 ( .A(n442), .ZN(y[1]) );
  AOI22_X1 U68 ( .A1(a[1]), .A2(n387), .B1(b[1]), .B2(n394), .ZN(n442) );
  INV_X1 U69 ( .A(n458), .ZN(y[5]) );
  AOI22_X1 U70 ( .A1(a[5]), .A2(n386), .B1(b[5]), .B2(n390), .ZN(n458) );
  INV_X1 U71 ( .A(n453), .ZN(y[2]) );
  AOI22_X1 U72 ( .A1(a[2]), .A2(n388), .B1(b[2]), .B2(n391), .ZN(n453) );
  INV_X1 U73 ( .A(n456), .ZN(y[3]) );
  AOI22_X1 U74 ( .A1(a[3]), .A2(sel), .B1(b[3]), .B2(n390), .ZN(n456) );
  INV_X1 U75 ( .A(n457), .ZN(y[4]) );
  AOI22_X1 U76 ( .A1(a[4]), .A2(n386), .B1(b[4]), .B2(n390), .ZN(n457) );
  BUF_X1 U77 ( .A(sel), .Z(n386) );
endmodule


module SHIFTER_M32_N5_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \temp_int_SH[4] , \SHMAG[5] , \MR_int[1][31] , \MR_int[1][30] ,
         \MR_int[1][29] , \MR_int[1][28] , \MR_int[1][27] , \MR_int[1][26] ,
         \MR_int[1][25] , \MR_int[1][24] , \MR_int[1][22] , \MR_int[1][21] ,
         \MR_int[1][16] , \MR_int[1][15] , \MR_int[1][14] , \MR_int[1][13] ,
         \MR_int[1][12] , \MR_int[1][11] , \MR_int[1][10] , \MR_int[1][9] ,
         \MR_int[1][8] , \MR_int[1][7] , \MR_int[1][6] , \MR_int[1][5] ,
         \MR_int[1][4] , \MR_int[1][3] , \MR_int[1][2] , \MR_int[1][1] ,
         \MR_int[2][31] , \MR_int[2][30] , \MR_int[2][29] , \MR_int[2][27] ,
         \MR_int[2][26] , \MR_int[2][25] , \MR_int[2][24] , \MR_int[2][23] ,
         \MR_int[2][22] , \MR_int[2][21] , \MR_int[2][20] , \MR_int[2][19] ,
         \MR_int[2][16] , \MR_int[2][15] , \MR_int[2][11] , \MR_int[2][10] ,
         \MR_int[2][9] , \MR_int[2][8] , \MR_int[2][7] , \MR_int[2][6] ,
         \MR_int[2][5] , \MR_int[2][4] , \MR_int[2][3] , \MR_int[2][2] ,
         \MR_int[2][1] , \MR_int[3][31] , \MR_int[3][30] , \MR_int[3][29] ,
         \MR_int[3][27] , \MR_int[3][26] , \MR_int[3][25] , \MR_int[3][24] ,
         \MR_int[3][23] , \MR_int[3][21] , \MR_int[3][20] , \MR_int[3][19] ,
         \MR_int[3][18] , \MR_int[3][17] , \MR_int[3][16] , \MR_int[3][15] ,
         \MR_int[3][12] , \MR_int[3][11] , \MR_int[3][10] , \MR_int[3][9] ,
         \MR_int[3][8] , \MR_int[3][7] , \MR_int[3][6] , \MR_int[3][4] ,
         \MR_int[3][3] , \MR_int[3][2] , \MR_int[3][1] , \MR_int[4][31] ,
         \MR_int[4][29] , \MR_int[4][28] , \MR_int[4][25] , \MR_int[4][24] ,
         \MR_int[4][22] , \MR_int[4][20] , \MR_int[4][19] , \MR_int[4][18] ,
         \MR_int[4][13] , \MR_int[4][12] , \MR_int[4][11] , \MR_int[4][10] ,
         \MR_int[4][8] , \MR_int[4][6] , \MR_int[4][4] , \MR_int[4][3] ,
         \MR_int[4][2] , \MR_int[5][3] , \MR_int[7][30] , \MR_int[7][29] ,
         \MR_int[7][24] , \MR_int[7][22] , \MR_int[7][20] , \MR_int[7][16] ,
         \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] , \ML_int[1][23] ,
         \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][19] , \ML_int[1][18] ,
         \ML_int[1][17] , \ML_int[1][16] , \ML_int[1][15] , \ML_int[1][14] ,
         \ML_int[1][13] , \ML_int[1][12] , \ML_int[1][11] , \ML_int[1][10] ,
         \ML_int[1][9] , \ML_int[1][8] , \ML_int[1][7] , \ML_int[1][6] ,
         \ML_int[1][5] , \ML_int[1][4] , \ML_int[1][3] , \ML_int[1][2] ,
         \ML_int[1][1] , \ML_int[1][0] , \ML_int[2][31] , \ML_int[2][30] ,
         \ML_int[2][29] , \ML_int[2][28] , \ML_int[2][26] , \ML_int[2][25] ,
         \ML_int[2][24] , \ML_int[2][23] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][17] , \ML_int[2][16] , \ML_int[2][15] ,
         \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] , \ML_int[2][11] ,
         \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] ,
         \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] ,
         \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] , \ML_int[3][31] ,
         \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] , \ML_int[3][27] ,
         \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] , \ML_int[3][23] ,
         \ML_int[3][21] , \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] ,
         \ML_int[3][16] , \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][15] ,
         \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] , \ML_int[4][11] ,
         \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] , \ML_int[5][31] ,
         \ML_int[5][30] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][18] , \ML_int[5][17] , \ML_int[7][29] , \ML_int[7][28] ,
         \ML_int[7][16] , \ML_int[7][14] , \ML_int[7][10] , \ML_int[7][9] ,
         \ML_int[7][7] , \ML_int[7][6] , \ML_int[7][5] , \ML_int[7][3] ,
         \ML_int[7][2] , \ML_int[7][1] , \ML_int[7][0] , n15, n80, n81, n82,
         n84, n85, n86, n87, n88, n90, n92, n98, n104, net60450, net60477,
         net60578, net60604, net60660, net60751, net60750, net60763, net60869,
         net60893, net61039, net61046, net61053, net61132, net61266, net61331,
         net61353, net61364, net61363, net61624, net61724, net61755, net61774,
         net61783, net61782, net61842, net61851, \ML_int[1][20] ,
         \ML_int[3][22] , \ML_int[2][22] , \ML_int[2][18] , net65464, net65465,
         \temp_int_SH[0] , net61465, n99, n97, n91, n101, n100,
         \MR_int[2][14] , \MR_int[4][30] , \MR_int[1][20] , \MR_int[1][18] ,
         net60718, \ML_int[7][13] , net61436, net60589, net60588,
         \MR_int[4][14] , \MR_int[3][22] , \MR_int[3][14] , \MR_int[2][18] ,
         n121, n122, n124, n125, n131, n132, n135, n136, n138, n139, n141,
         n142, n144, n145, n147, n148, n150, n151, n153, n154, n155, n156,
         n157, n158, n160, n161, n162, n163, n164, n168, n170, n171, n173,
         n174, n175, n178, n180, n181, n182, n183, n184, n186, n189, n192,
         n193, n195, n196, n197, n199, n200, n201, n204, n205, n207, n208,
         n211, n212, n213, n214, n215, n219, n220, n221, n223, n224, n225,
         n227, n228, n232, n233, n234, n235, n236, n237, n241, n243, n244,
         n245, n246, n250, n251, n252, n253, n255, n256, n257, n261, n264,
         n267, n270, n271, n272, n273, n274, n279, n282, n283, n284, n285,
         n286, n295, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n318,
         n319, n320, n321, n324, n325, n326, n327, n328, n329, n331, n332,
         n333, n334, n335, n336, n337, n338, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n369, n370, n375, n376, n377, n378, n379, n380, n381, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n403, n404, n405, n406, n407,
         n409, n410, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n502, n503, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n532, n535, n536, n537, n538,
         n539, n540, n542, n543, n544, n545, n546, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n565, n566, n567, n568, n569, n570, n571, n572, n574, n575, n576,
         n577, n578, n579, n580, n581, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n611, n622,
         n623, n624, n627, n628, net135734, net141444, net141501, net141507,
         net141562, net141573, n290, n289, n288, n287, n109, n108, n107, n106,
         n96, n89, \MR_int[1][19] , net60313, n292, n291, n110,
         \temp_int_SH[3] , \temp_int_SH[1] , net60576, n95, \MR_int[1][17] ,
         \temp_int_SH[2] , n548, n547, n260, \MR_int[2][17] , \MR_int[2][13] ,
         n83, n340, \ML_int[7][4] , \MR_int[3][13] , n128, n127,
         \MR_int[4][5] , \MR_int[3][5] , n656, n660, n661, n662, n664, n666,
         n667, n668, n669, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n684, n686, n688, n689, n690, n691, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n706, n707, n708, n709, n712, n713,
         n714, n715, n717, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n743, n744, n745, n759, n760, n761, n762, n763, n800, n801,
         n802, n803, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051;

  MUX2_X1 M1_3_3 ( .A(\MR_int[3][3] ), .B(\MR_int[3][11] ), .S(n1009), .Z(
        \MR_int[4][3] ) );
  MUX2_X1 M1_3_2 ( .A(\MR_int[3][2] ), .B(\MR_int[3][10] ), .S(n1007), .Z(
        \MR_int[4][2] ) );
  MUX2_X1 M1_2_6_0 ( .A(\MR_int[2][6] ), .B(\MR_int[2][10] ), .S(n969), .Z(
        \MR_int[3][6] ) );
  MUX2_X1 M1_2_4_0 ( .A(\MR_int[2][4] ), .B(\MR_int[2][8] ), .S(n969), .Z(
        \MR_int[3][4] ) );
  MUX2_X1 M1_2_3 ( .A(\MR_int[2][3] ), .B(\MR_int[2][7] ), .S(n969), .Z(
        \MR_int[3][3] ) );
  MUX2_X1 M1_1_11_0 ( .A(\MR_int[1][11] ), .B(\MR_int[1][13] ), .S(n988), .Z(
        \MR_int[2][11] ) );
  MUX2_X1 M1_1_10_0 ( .A(\MR_int[1][10] ), .B(\MR_int[1][12] ), .S(n988), .Z(
        \MR_int[2][10] ) );
  MUX2_X1 M1_1_4_0 ( .A(\MR_int[1][4] ), .B(\MR_int[1][6] ), .S(n988), .Z(
        \MR_int[2][4] ) );
  MUX2_X1 M1_1_3_0 ( .A(\MR_int[1][3] ), .B(\MR_int[1][5] ), .S(n988), .Z(
        \MR_int[2][3] ) );
  MUX2_X1 M1_1_1 ( .A(\MR_int[1][1] ), .B(\ML_int[1][4] ), .S(n988), .Z(
        \MR_int[2][1] ) );
  MUX2_X1 M1_0_29_0 ( .A(A[29]), .B(A[30]), .S(n1032), .Z(\MR_int[1][29] ) );
  MUX2_X1 M1_0_28_0 ( .A(A[28]), .B(A[29]), .S(n1032), .Z(\MR_int[1][28] ) );
  MUX2_X1 M1_0_24_0 ( .A(A[24]), .B(A[25]), .S(n1032), .Z(\MR_int[1][24] ) );
  MUX2_X1 M1_0_22_0 ( .A(A[22]), .B(A[23]), .S(net141501), .Z(\MR_int[1][22] )
         );
  MUX2_X1 M1_0_9_0 ( .A(A[9]), .B(A[10]), .S(n1045), .Z(\MR_int[1][9] ) );
  MUX2_X1 M1_0_8_0 ( .A(A[8]), .B(A[9]), .S(n1045), .Z(\MR_int[1][8] ) );
  MUX2_X1 M1_0_6_0 ( .A(A[6]), .B(A[7]), .S(n1032), .Z(\MR_int[1][6] ) );
  MUX2_X1 M1_0_5_0 ( .A(A[5]), .B(A[6]), .S(n1032), .Z(\MR_int[1][5] ) );
  MUX2_X1 M1_0_4_0 ( .A(A[4]), .B(A[5]), .S(n1032), .Z(\MR_int[1][4] ) );
  MUX2_X1 M1_0_2_0 ( .A(A[2]), .B(A[3]), .S(net141501), .Z(\MR_int[1][2] ) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n1017), .Z(
        \ML_int[5][25] ) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(n1028), .S(n1017), .Z(
        \ML_int[5][18] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n998), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n981), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n980), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(n297), .S(n980), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n981), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(net135734), .Z(\ML_int[1][31] )
         );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(net135734), .Z(\ML_int[1][29] )
         );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n1039), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n1039), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n1039), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(net61851), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(net61851), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(net135734), .Z(\ML_int[1][16] )
         );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(net135734), .Z(\ML_int[1][15] )
         );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n1039), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(\temp_int_SH[0] ), .Z(
        \ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(net135734), .Z(\ML_int[1][12] )
         );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(\temp_int_SH[0] ), .Z(
        \ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(net61851), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n1039), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(net135734), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(\temp_int_SH[0] ), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(\temp_int_SH[0] ), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(net61851), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n1039), .Z(\ML_int[1][1] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n1039), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n1039), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n1039), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n981), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n729), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_13_0 ( .A(A[13]), .B(A[14]), .S(n1045), .Z(\MR_int[1][13] ) );
  MUX2_X1 M1_0_1_0 ( .A(A[1]), .B(A[2]), .S(n1032), .Z(\MR_int[1][1] ) );
  MUX2_X1 M1_3_22_0 ( .A(n727), .B(\MR_int[3][30] ), .S(n1009), .Z(
        \MR_int[4][22] ) );
  MUX2_X1 M1_3_11_0 ( .A(\MR_int[3][11] ), .B(\MR_int[3][19] ), .S(n1009), .Z(
        \MR_int[4][11] ) );
  MUX2_X1 M1_3_14_0 ( .A(n669), .B(n727), .S(n1008), .Z(\MR_int[4][14] ) );
  MUX2_X1 M1_2_27_0 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n969), .Z(
        \MR_int[3][27] ) );
  MUX2_X1 U3 ( .A(\ML_int[2][26] ), .B(\ML_int[2][30] ), .S(n969), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 U9 ( .A(\MR_int[2][6] ), .B(\MR_int[2][2] ), .S(n959), .Z(
        \MR_int[3][2] ) );
  MUX2_X1 U47 ( .A(\ML_int[3][23] ), .B(\ML_int[3][31] ), .S(n1009), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 U78 ( .A(\ML_int[7][16] ), .B(\MR_int[7][16] ), .S(SH[31]), .Z(B[16]) );
  MUX2_X1 U93 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n998), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 U127 ( .A(A[22]), .B(A[23]), .S(net141501), .Z(n186) );
  MUX2_X1 U197 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n969), .Z(n236)
         );
  MUX2_X1 U204 ( .A(\MR_int[3][10] ), .B(\MR_int[3][18] ), .S(n1009), .Z(
        \MR_int[4][10] ) );
  MUX2_X1 U226 ( .A(\MR_int[2][11] ), .B(\MR_int[2][7] ), .S(n959), .Z(
        \MR_int[3][7] ) );
  MUX2_X1 U228 ( .A(\MR_int[1][9] ), .B(\MR_int[1][7] ), .S(n981), .Z(
        \MR_int[2][7] ) );
  MUX2_X1 U235 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n980), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 U236 ( .A(\ML_int[2][18] ), .B(\ML_int[2][22] ), .S(n969), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 U241 ( .A(\ML_int[1][11] ), .B(n728), .S(n988), .Z(n264) );
  MUX2_X1 U248 ( .A(\ML_int[3][9] ), .B(\ML_int[3][17] ), .S(n1008), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 U254 ( .A(\ML_int[1][24] ), .B(\ML_int[1][26] ), .S(n988), .Z(
        \ML_int[2][26] ) );
  NAND3_X1 U269 ( .A1(\ML_int[5][25] ), .A2(n85), .A3(n948), .ZN(n336) );
  NAND3_X1 U271 ( .A1(\ML_int[5][24] ), .A2(n85), .A3(n948), .ZN(n527) );
  MUX2_X1 U288 ( .A(\MR_int[1][20] ), .B(\MR_int[1][18] ), .S(n981), .Z(
        \MR_int[2][18] ) );
  MUX2_X1 U294 ( .A(\MR_int[3][22] ), .B(\MR_int[3][30] ), .S(n1007), .Z(
        net61774) );
  MUX2_X1 U370 ( .A(\MR_int[3][4] ), .B(\MR_int[3][12] ), .S(n1009), .Z(
        \MR_int[4][4] ) );
  MUX2_X1 U374 ( .A(A[26]), .B(A[25]), .S(net135734), .Z(n297) );
  MUX2_X1 U389 ( .A(A[11]), .B(A[10]), .S(net135734), .Z(\MR_int[1][10] ) );
  MUX2_X1 U448 ( .A(A[8]), .B(A[7]), .S(n1039), .Z(\MR_int[1][7] ) );
  MUX2_X1 U493 ( .A(A[28]), .B(A[27]), .S(net135734), .Z(\MR_int[1][27] ) );
  MUX2_X1 U557 ( .A(A[4]), .B(A[3]), .S(net135734), .Z(\MR_int[1][3] ) );
  MUX2_X1 U558 ( .A(A[30]), .B(A[31]), .S(n1032), .Z(\MR_int[1][30] ) );
  MUX2_X1 U565 ( .A(A[13]), .B(A[12]), .S(n1039), .Z(\MR_int[1][12] ) );
  MUX2_X1 U601 ( .A(\MR_int[1][12] ), .B(\MR_int[1][14] ), .S(n988), .Z(n410)
         );
  MUX2_X1 U621 ( .A(A[27]), .B(A[26]), .S(n1039), .Z(n424) );
  MUX2_X1 U734 ( .A(A[16]), .B(A[15]), .S(n729), .Z(\MR_int[1][15] ) );
  MUX2_X1 U768 ( .A(A[15]), .B(A[14]), .S(n729), .Z(\MR_int[1][14] ) );
  MUX2_X1 U777 ( .A(\MR_int[3][16] ), .B(\MR_int[3][8] ), .S(n998), .Z(
        \MR_int[4][8] ) );
  MUX2_X1 U913 ( .A(A[23]), .B(A[24]), .S(n1045), .Z(n601) );
  MUX2_X1 U299 ( .A(n424), .B(\ML_int[1][25] ), .S(n980), .Z(n250) );
  MUX2_X1 U732 ( .A(\ML_int[7][29] ), .B(\MR_int[7][29] ), .S(SH[31]), .Z(
        B[29]) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n959), .Z(
        \ML_int[3][4] ) );
  NAND3_X1 U365 ( .A1(SH[16]), .A2(SH[15]), .A3(SH[14]), .ZN(net60751) );
  NAND3_X1 U364 ( .A1(SH[18]), .A2(SH[17]), .A3(SH[19]), .ZN(net61363) );
  NAND3_X1 U281 ( .A1(SH[22]), .A2(SH[21]), .A3(SH[20]), .ZN(net61364) );
  MUX2_X1 M1_0_20_0 ( .A(A[20]), .B(A[21]), .S(n1032), .Z(\MR_int[1][20] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(net61851), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(net135734), .Z(\ML_int[1][21] )
         );
  NAND3_X1 U367 ( .A1(SH[8]), .A2(SH[7]), .A3(SH[9]), .ZN(net65464) );
  NAND3_X1 U368 ( .A1(SH[30]), .A2(SH[29]), .A3(SH[6]), .ZN(net65465) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(net61851), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n1039), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16_0 ( .A(A[16]), .B(A[17]), .S(n1032), .Z(\MR_int[1][16] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(\temp_int_SH[0] ), .Z(
        \ML_int[1][18] ) );
  MUX2_X1 M1_0_25_0 ( .A(A[25]), .B(A[26]), .S(n1032), .Z(\MR_int[1][25] ) );
  MUX2_X1 M1_0_17_0 ( .A(A[17]), .B(A[18]), .S(n1032), .Z(\MR_int[1][17] ) );
  MUX2_X1 M1_2_5_0 ( .A(\MR_int[2][5] ), .B(\MR_int[2][9] ), .S(n969), .Z(
        \MR_int[3][5] ) );
  MUX2_X1 U29 ( .A(A[30]), .B(A[29]), .S(\temp_int_SH[0] ), .Z(\ML_int[1][30] ) );
  MUX2_X1 U42 ( .A(\MR_int[3][12] ), .B(\MR_int[3][20] ), .S(n1009), .Z(
        \MR_int[4][12] ) );
  MUX2_X1 U44 ( .A(\MR_int[1][13] ), .B(\MR_int[1][15] ), .S(n988), .Z(
        \MR_int[2][13] ) );
  MUX2_X1 U46 ( .A(A[19]), .B(A[18]), .S(\temp_int_SH[0] ), .Z(\MR_int[1][18] ) );
  NAND3_X1 U61 ( .A1(n422), .A2(n225), .A3(n423), .ZN(n163) );
  MUX2_X1 U67 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n959), .Z(
        \ML_int[3][26] ) );
  NAND3_X1 U74 ( .A1(n232), .A2(n233), .A3(n594), .ZN(B[9]) );
  NAND3_X1 U81 ( .A1(n363), .A2(n409), .A3(n364), .ZN(\ML_int[4][9] ) );
  MUX2_X1 U96 ( .A(\MR_int[1][20] ), .B(\MR_int[1][18] ), .S(n981), .Z(
        net61353) );
  MUX2_X1 U154 ( .A(\MR_int[2][17] ), .B(\MR_int[2][13] ), .S(n959), .Z(
        \MR_int[3][13] ) );
  MUX2_X1 U169 ( .A(\MR_int[2][13] ), .B(\MR_int[2][17] ), .S(n969), .Z(
        net141562) );
  MUX2_X1 U199 ( .A(A[20]), .B(A[19]), .S(n1039), .Z(\MR_int[1][19] ) );
  MUX2_X1 U217 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n959), .Z(
        net141573) );
  MUX2_X1 U221 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n969), .Z(n725)
         );
  MUX2_X1 U222 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n969), .Z(n726)
         );
  MUX2_X1 U225 ( .A(A[13]), .B(A[12]), .S(\temp_int_SH[0] ), .Z(n728) );
  MUX2_X1 U227 ( .A(A[27]), .B(A[26]), .S(n1039), .Z(\MR_int[1][26] ) );
  MUX2_X1 U243 ( .A(A[12]), .B(A[11]), .S(n1039), .Z(\MR_int[1][11] ) );
  MUX2_X1 U244 ( .A(A[28]), .B(A[29]), .S(net141501), .Z(n732) );
  MUX2_X1 U582 ( .A(\MR_int[1][11] ), .B(\MR_int[1][9] ), .S(n980), .Z(
        \MR_int[2][9] ) );
  MUX2_X1 U608 ( .A(A[22]), .B(A[21]), .S(net135734), .Z(\MR_int[1][21] ) );
  MUX2_X1 U337 ( .A(\MR_int[2][30] ), .B(\MR_int[2][26] ), .S(n959), .Z(
        \MR_int[3][26] ) );
  AND2_X1 U4 ( .A1(net61465), .A2(n92), .ZN(\SHMAG[5] ) );
  AND2_X1 U5 ( .A1(n967), .A2(n1008), .ZN(n365) );
  INV_X1 U6 ( .A(n960), .ZN(n967) );
  INV_X1 U7 ( .A(n999), .ZN(n1007) );
  INV_X1 U8 ( .A(n999), .ZN(n1008) );
  INV_X1 U10 ( .A(n960), .ZN(n969) );
  INV_X1 U11 ( .A(n960), .ZN(n968) );
  INV_X1 U12 ( .A(n999), .ZN(n1009) );
  NAND2_X1 U13 ( .A1(\MR_int[3][31] ), .A2(n1007), .ZN(n603) );
  NAND2_X1 U14 ( .A1(n730), .A2(n1008), .ZN(n628) );
  NAND2_X1 U15 ( .A1(\MR_int[3][23] ), .A2(n184), .ZN(n182) );
  AND2_X1 U16 ( .A1(n1000), .A2(n1014), .ZN(n184) );
  AND2_X1 U17 ( .A1(n960), .A2(n1008), .ZN(n357) );
  AND2_X1 U18 ( .A1(n1000), .A2(n1014), .ZN(n175) );
  AND2_X1 U19 ( .A1(n986), .A2(n969), .ZN(n731) );
  AND2_X1 U20 ( .A1(n1000), .A2(n155), .ZN(\MR_int[4][30] ) );
  INV_X1 U21 ( .A(n88), .ZN(n1030) );
  INV_X1 U22 ( .A(n87), .ZN(n1038) );
  INV_X1 U23 ( .A(n81), .ZN(n1029) );
  INV_X1 U24 ( .A(n84), .ZN(n1034) );
  OR2_X1 U25 ( .A1(n1014), .A2(n491), .ZN(n245) );
  INV_X1 U26 ( .A(n982), .ZN(n987) );
  INV_X1 U27 ( .A(n982), .ZN(n986) );
  INV_X1 U28 ( .A(n982), .ZN(n988) );
  BUF_X1 U30 ( .A(n1010), .Z(n1012) );
  BUF_X1 U31 ( .A(n1010), .Z(n1013) );
  BUF_X1 U32 ( .A(n1011), .Z(n1014) );
  NOR2_X1 U33 ( .A1(n968), .A2(n1027), .ZN(n155) );
  AOI21_X1 U34 ( .B1(n468), .B2(n467), .A(n1014), .ZN(n690) );
  NAND2_X1 U35 ( .A1(\MR_int[3][9] ), .A2(n990), .ZN(n467) );
  OAI21_X1 U36 ( .B1(n1040), .B2(n689), .A(n1009), .ZN(n468) );
  INV_X1 U37 ( .A(n565), .ZN(n1040) );
  NOR2_X1 U38 ( .A1(n969), .A2(n392), .ZN(\MR_int[3][31] ) );
  BUF_X1 U39 ( .A(n1001), .Z(n999) );
  BUF_X1 U40 ( .A(n961), .Z(n960) );
  NOR2_X1 U41 ( .A1(n325), .A2(n84), .ZN(\ML_int[7][3] ) );
  NOR2_X1 U43 ( .A1(n80), .A2(n325), .ZN(\ML_int[7][7] ) );
  BUF_X1 U45 ( .A(n961), .Z(n959) );
  NOR2_X1 U48 ( .A1(n1042), .A2(n1017), .ZN(n733) );
  NAND2_X1 U49 ( .A1(\ML_int[3][0] ), .A2(n1007), .ZN(n88) );
  NAND2_X1 U50 ( .A1(\ML_int[3][1] ), .A2(n1007), .ZN(n87) );
  NAND2_X1 U51 ( .A1(\ML_int[3][6] ), .A2(n1007), .ZN(n81) );
  NAND2_X1 U52 ( .A1(\ML_int[3][3] ), .A2(n1007), .ZN(n84) );
  NAND2_X1 U53 ( .A1(\ML_int[3][2] ), .A2(n1007), .ZN(n86) );
  NAND2_X1 U54 ( .A1(\ML_int[3][5] ), .A2(n1007), .ZN(n82) );
  NOR2_X1 U55 ( .A1(n969), .A2(n1027), .ZN(\MR_int[3][30] ) );
  BUF_X1 U56 ( .A(n964), .Z(n950) );
  BUF_X1 U57 ( .A(n963), .Z(n953) );
  BUF_X1 U58 ( .A(n963), .Z(n952) );
  BUF_X1 U59 ( .A(n964), .Z(n951) );
  BUF_X1 U60 ( .A(n964), .Z(n949) );
  BUF_X1 U62 ( .A(n962), .Z(n955) );
  BUF_X1 U63 ( .A(n962), .Z(n957) );
  BUF_X1 U64 ( .A(n963), .Z(n954) );
  BUF_X1 U65 ( .A(n962), .Z(n956) );
  BUF_X1 U66 ( .A(n1004), .Z(n991) );
  BUF_X1 U68 ( .A(n1004), .Z(n989) );
  BUF_X1 U69 ( .A(n1004), .Z(n990) );
  BUF_X1 U70 ( .A(n1003), .Z(n993) );
  BUF_X1 U71 ( .A(n1003), .Z(n994) );
  BUF_X1 U72 ( .A(n1002), .Z(n996) );
  BUF_X1 U73 ( .A(n1003), .Z(n992) );
  BUF_X1 U75 ( .A(n1002), .Z(n995) );
  BUF_X1 U76 ( .A(n961), .Z(n958) );
  BUF_X1 U77 ( .A(n1002), .Z(n997) );
  BUF_X1 U79 ( .A(n1001), .Z(n1000) );
  BUF_X1 U80 ( .A(n1001), .Z(n998) );
  NAND2_X1 U82 ( .A1(n345), .A2(n365), .ZN(n363) );
  OR2_X1 U83 ( .A1(n466), .A2(n1000), .ZN(n364) );
  NAND2_X1 U84 ( .A1(\ML_int[3][1] ), .A2(n993), .ZN(n409) );
  NAND2_X1 U85 ( .A1(\ML_int[3][7] ), .A2(n1007), .ZN(n80) );
  NAND2_X1 U86 ( .A1(\MR_int[3][19] ), .A2(n989), .ZN(n604) );
  BUF_X1 U87 ( .A(n1011), .Z(n1015) );
  NAND2_X1 U88 ( .A1(n445), .A2(n444), .ZN(\MR_int[3][23] ) );
  NAND2_X1 U89 ( .A1(n1023), .A2(n565), .ZN(\MR_int[3][17] ) );
  INV_X1 U90 ( .A(n689), .ZN(n1023) );
  NAND2_X1 U91 ( .A1(n484), .A2(n485), .ZN(n730) );
  NAND2_X1 U92 ( .A1(n437), .A2(n438), .ZN(\ML_int[4][11] ) );
  NAND2_X1 U94 ( .A1(\ML_int[3][3] ), .A2(n993), .ZN(n438) );
  NAND2_X1 U95 ( .A1(\ML_int[3][11] ), .A2(n1009), .ZN(n437) );
  NAND2_X1 U97 ( .A1(n345), .A2(n968), .ZN(n465) );
  NAND2_X1 U98 ( .A1(\ML_int[3][0] ), .A2(n990), .ZN(n491) );
  NAND2_X1 U99 ( .A1(\ML_int[3][18] ), .A2(n1007), .ZN(n369) );
  NAND2_X1 U100 ( .A1(\ML_int[3][19] ), .A2(n1007), .ZN(n425) );
  NAND2_X1 U101 ( .A1(n551), .A2(n550), .ZN(\ML_int[4][14] ) );
  NAND2_X1 U102 ( .A1(\ML_int[3][6] ), .A2(n994), .ZN(n551) );
  NAND2_X1 U103 ( .A1(\ML_int[3][14] ), .A2(n1009), .ZN(n550) );
  NAND2_X1 U104 ( .A1(net61132), .A2(n475), .ZN(\ML_int[4][15] ) );
  NAND2_X1 U105 ( .A1(\ML_int[3][7] ), .A2(n995), .ZN(n475) );
  NAND2_X1 U106 ( .A1(\ML_int[3][15] ), .A2(n1008), .ZN(net61132) );
  NAND2_X1 U107 ( .A1(n138), .A2(n139), .ZN(\ML_int[4][10] ) );
  NAND2_X1 U108 ( .A1(\ML_int[3][2] ), .A2(n994), .ZN(n139) );
  NAND2_X1 U109 ( .A1(\ML_int[3][10] ), .A2(n1009), .ZN(n138) );
  NAND2_X1 U110 ( .A1(n174), .A2(n1009), .ZN(n423) );
  NAND2_X1 U111 ( .A1(n445), .A2(n444), .ZN(n174) );
  NAND2_X1 U112 ( .A1(\MR_int[3][21] ), .A2(n990), .ZN(n606) );
  NAND2_X1 U113 ( .A1(\ML_int[4][11] ), .A2(n1016), .ZN(n701) );
  NAND2_X1 U114 ( .A1(\ML_int[3][10] ), .A2(n991), .ZN(n370) );
  NAND2_X1 U115 ( .A1(\ML_int[3][11] ), .A2(n992), .ZN(n426) );
  NAND2_X1 U116 ( .A1(n1033), .A2(n1016), .ZN(n125) );
  INV_X1 U117 ( .A(n82), .ZN(n1033) );
  NAND2_X1 U118 ( .A1(\ML_int[4][14] ), .A2(n1016), .ZN(n715) );
  NAND2_X1 U119 ( .A1(\ML_int[5][22] ), .A2(n493), .ZN(n495) );
  NAND2_X1 U120 ( .A1(n697), .A2(n698), .ZN(\ML_int[5][22] ) );
  NAND2_X1 U121 ( .A1(\ML_int[4][22] ), .A2(n1012), .ZN(n697) );
  NAND2_X1 U122 ( .A1(n1029), .A2(n1016), .ZN(n698) );
  NAND2_X1 U123 ( .A1(n400), .A2(n399), .ZN(\ML_int[4][20] ) );
  NAND2_X1 U124 ( .A1(n251), .A2(n996), .ZN(n400) );
  NAND2_X1 U125 ( .A1(n253), .A2(n1007), .ZN(n399) );
  NAND2_X1 U126 ( .A1(n430), .A2(n429), .ZN(\ML_int[4][27] ) );
  NAND2_X1 U128 ( .A1(\ML_int[3][19] ), .A2(n997), .ZN(n429) );
  NAND2_X1 U129 ( .A1(\ML_int[3][27] ), .A2(n1008), .ZN(n430) );
  NAND2_X1 U130 ( .A1(n480), .A2(n481), .ZN(\ML_int[3][27] ) );
  NAND2_X1 U131 ( .A1(\ML_int[5][17] ), .A2(n379), .ZN(n450) );
  NAND2_X1 U132 ( .A1(n360), .A2(n361), .ZN(\ML_int[5][17] ) );
  NAND2_X1 U133 ( .A1(\ML_int[4][17] ), .A2(n1013), .ZN(n360) );
  NAND2_X1 U134 ( .A1(n1038), .A2(n1016), .ZN(n361) );
  NAND2_X1 U135 ( .A1(\ML_int[5][18] ), .A2(n227), .ZN(n436) );
  INV_X1 U136 ( .A(n86), .ZN(n1028) );
  NAND2_X1 U137 ( .A1(n369), .A2(n370), .ZN(\ML_int[4][18] ) );
  NAND2_X1 U138 ( .A1(\ML_int[5][20] ), .A2(n227), .ZN(n443) );
  NAND2_X1 U139 ( .A1(n366), .A2(n367), .ZN(\ML_int[5][20] ) );
  NAND2_X1 U140 ( .A1(\ML_int[4][20] ), .A2(n1013), .ZN(n366) );
  NAND2_X1 U141 ( .A1(n309), .A2(n1016), .ZN(n367) );
  NAND2_X1 U142 ( .A1(\ML_int[5][23] ), .A2(n379), .ZN(n514) );
  NAND2_X1 U143 ( .A1(n471), .A2(n472), .ZN(\ML_int[5][23] ) );
  OR2_X1 U144 ( .A1(n80), .A2(n1015), .ZN(n472) );
  NAND2_X1 U145 ( .A1(\ML_int[4][23] ), .A2(n1012), .ZN(n471) );
  NAND2_X1 U146 ( .A1(n513), .A2(n512), .ZN(\ML_int[4][23] ) );
  NAND2_X1 U147 ( .A1(\ML_int[3][15] ), .A2(n995), .ZN(n512) );
  NAND2_X1 U148 ( .A1(\ML_int[3][23] ), .A2(n1008), .ZN(n513) );
  NAND2_X1 U149 ( .A1(n431), .A2(n432), .ZN(\ML_int[4][24] ) );
  NAND2_X1 U150 ( .A1(\ML_int[3][16] ), .A2(n996), .ZN(n432) );
  NAND2_X1 U151 ( .A1(\ML_int[3][24] ), .A2(n1008), .ZN(n431) );
  NAND2_X1 U152 ( .A1(n341), .A2(n342), .ZN(\ML_int[3][24] ) );
  AND2_X1 U153 ( .A1(n1008), .A2(n1017), .ZN(n745) );
  OR2_X1 U155 ( .A1(n1017), .A2(n603), .ZN(n183) );
  NAND2_X1 U156 ( .A1(\MR_int[4][28] ), .A2(n1012), .ZN(n592) );
  NAND2_X1 U157 ( .A1(\MR_int[4][29] ), .A2(n1012), .ZN(n456) );
  NAND2_X1 U158 ( .A1(\MR_int[3][15] ), .A2(n993), .ZN(n422) );
  AND2_X1 U159 ( .A1(n1000), .A2(n205), .ZN(n664) );
  AND2_X1 U160 ( .A1(n622), .A2(\ML_int[4][13] ), .ZN(\ML_int[7][13] ) );
  AND2_X1 U161 ( .A1(net141573), .A2(n1007), .ZN(n309) );
  AND2_X1 U162 ( .A1(\ML_int[3][16] ), .A2(n158), .ZN(n161) );
  AND2_X1 U163 ( .A1(n1009), .A2(n252), .ZN(n158) );
  AND2_X1 U164 ( .A1(\ML_int[3][8] ), .A2(n199), .ZN(n160) );
  AND2_X1 U165 ( .A1(n1000), .A2(n252), .ZN(n199) );
  AND2_X1 U166 ( .A1(n606), .A2(n607), .ZN(n675) );
  AND2_X1 U167 ( .A1(n303), .A2(n304), .ZN(n674) );
  NAND2_X1 U168 ( .A1(\ML_int[4][19] ), .A2(n1012), .ZN(n303) );
  NAND2_X1 U170 ( .A1(n1034), .A2(n1016), .ZN(n304) );
  NAND2_X1 U171 ( .A1(n425), .A2(n426), .ZN(\ML_int[4][19] ) );
  NAND2_X1 U172 ( .A1(n484), .A2(n485), .ZN(\MR_int[3][24] ) );
  NAND2_X1 U173 ( .A1(\ML_int[3][8] ), .A2(n246), .ZN(n244) );
  AND2_X1 U174 ( .A1(n1007), .A2(n1017), .ZN(n246) );
  NAND2_X1 U175 ( .A1(n328), .A2(n329), .ZN(\ML_int[7][16] ) );
  OR2_X1 U176 ( .A1(n1042), .A2(n362), .ZN(n329) );
  NOR2_X1 U177 ( .A1(n160), .A2(n161), .ZN(n328) );
  NAND2_X1 U178 ( .A1(n1030), .A2(n1017), .ZN(n362) );
  NAND2_X1 U179 ( .A1(n661), .A2(n662), .ZN(\MR_int[7][16] ) );
  OR2_X1 U180 ( .A1(n1043), .A2(n243), .ZN(n662) );
  NAND2_X1 U181 ( .A1(\MR_int[3][17] ), .A2(n664), .ZN(n661) );
  INV_X1 U182 ( .A(n205), .ZN(n1043) );
  NAND2_X1 U183 ( .A1(n735), .A2(n734), .ZN(\ML_int[7][29] ) );
  NAND2_X1 U184 ( .A1(\ML_int[4][29] ), .A2(n733), .ZN(n735) );
  NAND2_X1 U185 ( .A1(\ML_int[4][13] ), .A2(n736), .ZN(n734) );
  NAND2_X1 U186 ( .A1(n386), .A2(n387), .ZN(\ML_int[4][29] ) );
  INV_X1 U187 ( .A(n686), .ZN(n1020) );
  AOI21_X1 U188 ( .B1(n702), .B2(n701), .A(n1021), .ZN(n686) );
  INV_X1 U189 ( .A(n493), .ZN(n1021) );
  NAND2_X1 U190 ( .A1(\ML_int[4][27] ), .A2(n1013), .ZN(n702) );
  INV_X1 U191 ( .A(net141501), .ZN(n1039) );
  INV_X1 U192 ( .A(\temp_int_SH[0] ), .ZN(n1032) );
  NAND2_X1 U193 ( .A1(n85), .A2(n1012), .ZN(n325) );
  OAI22_X1 U194 ( .A1(n1037), .A2(n671), .B1(net61039), .B2(n1009), .ZN(n688)
         );
  INV_X1 U195 ( .A(n348), .ZN(n1037) );
  NAND2_X1 U196 ( .A1(n969), .A2(n989), .ZN(n671) );
  AOI21_X1 U198 ( .B1(n547), .B2(n548), .A(n969), .ZN(n689) );
  BUF_X1 U200 ( .A(\temp_int_SH[4] ), .Z(n1017) );
  AND2_X1 U201 ( .A1(n85), .A2(n1014), .ZN(n622) );
  BUF_X1 U202 ( .A(\temp_int_SH[4] ), .Z(n1016) );
  OAI21_X1 U203 ( .B1(n969), .B2(n1036), .A(n503), .ZN(\ML_int[3][19] ) );
  INV_X1 U205 ( .A(\ML_int[2][15] ), .ZN(n1036) );
  NAND2_X1 U206 ( .A1(\ML_int[2][19] ), .A2(n968), .ZN(n503) );
  NAND2_X1 U207 ( .A1(n353), .A2(n352), .ZN(\ML_int[2][19] ) );
  AOI22_X1 U208 ( .A1(\MR_int[4][11] ), .A2(n383), .B1(n520), .B2(n261), .ZN(
        n584) );
  AND2_X1 U209 ( .A1(n1017), .A2(n405), .ZN(n383) );
  NOR2_X1 U210 ( .A1(n1009), .A2(n448), .ZN(n520) );
  OAI21_X1 U211 ( .B1(n219), .B2(n968), .A(n464), .ZN(\ML_int[3][23] ) );
  AND2_X1 U212 ( .A1(n352), .A2(n353), .ZN(n219) );
  NAND2_X1 U213 ( .A1(\ML_int[2][23] ), .A2(n969), .ZN(n464) );
  NOR2_X1 U214 ( .A1(n988), .A2(n1031), .ZN(\MR_int[2][31] ) );
  NAND2_X1 U215 ( .A1(n470), .A2(n469), .ZN(\ML_int[5][24] ) );
  AND2_X1 U216 ( .A1(n244), .A2(n245), .ZN(n469) );
  NAND2_X1 U218 ( .A1(\ML_int[4][24] ), .A2(n1012), .ZN(n470) );
  NAND2_X1 U219 ( .A1(n1035), .A2(n488), .ZN(\ML_int[4][25] ) );
  INV_X1 U220 ( .A(n688), .ZN(n1035) );
  AOI21_X1 U223 ( .B1(n193), .B2(n192), .A(n1014), .ZN(n684) );
  NAND2_X1 U224 ( .A1(\MR_int[3][7] ), .A2(n990), .ZN(n192) );
  NAND2_X1 U229 ( .A1(\MR_int[3][15] ), .A2(n1007), .ZN(n193) );
  NAND2_X1 U230 ( .A1(n200), .A2(n505), .ZN(n345) );
  AND2_X1 U231 ( .A1(n948), .A2(n85), .ZN(n493) );
  BUF_X1 U232 ( .A(n983), .Z(n982) );
  BUF_X1 U233 ( .A(n983), .Z(n981) );
  NAND2_X1 U234 ( .A1(\MR_int[2][27] ), .A2(n968), .ZN(n444) );
  NAND2_X1 U237 ( .A1(\MR_int[2][21] ), .A2(n968), .ZN(n565) );
  BUF_X1 U238 ( .A(n983), .Z(n980) );
  NAND2_X1 U239 ( .A1(n623), .A2(n967), .ZN(n484) );
  BUF_X1 U240 ( .A(n984), .Z(n974) );
  BUF_X1 U242 ( .A(n984), .Z(n975) );
  BUF_X1 U245 ( .A(n984), .Z(n973) );
  BUF_X1 U246 ( .A(n983), .Z(n978) );
  BUF_X1 U247 ( .A(n984), .Z(n977) );
  BUF_X1 U249 ( .A(n983), .Z(n979) );
  BUF_X1 U250 ( .A(n984), .Z(n976) );
  BUF_X1 U251 ( .A(n985), .Z(n972) );
  BUF_X1 U252 ( .A(n985), .Z(n971) );
  BUF_X1 U253 ( .A(n985), .Z(n970) );
  NAND2_X1 U255 ( .A1(n433), .A2(n434), .ZN(\ML_int[3][8] ) );
  NAND2_X1 U256 ( .A1(\ML_int[2][4] ), .A2(n952), .ZN(n434) );
  NAND2_X1 U257 ( .A1(\ML_int[2][8] ), .A2(n968), .ZN(n433) );
  NAND2_X1 U258 ( .A1(n85), .A2(n946), .ZN(n672) );
  INV_X1 U259 ( .A(n729), .ZN(n1045) );
  NAND2_X1 U260 ( .A1(\MR_int[2][24] ), .A2(n949), .ZN(n485) );
  NAND2_X1 U261 ( .A1(\MR_int[2][14] ), .A2(n949), .ZN(net60589) );
  NAND2_X1 U262 ( .A1(\MR_int[3][18] ), .A2(n989), .ZN(n575) );
  AND2_X1 U263 ( .A1(n1015), .A2(n85), .ZN(n252) );
  AND2_X1 U264 ( .A1(n85), .A2(n948), .ZN(n227) );
  AND2_X1 U265 ( .A1(n85), .A2(n948), .ZN(n379) );
  NAND2_X1 U266 ( .A1(\MR_int[2][23] ), .A2(n950), .ZN(n445) );
  NAND2_X1 U267 ( .A1(\MR_int[3][20] ), .A2(n989), .ZN(n522) );
  NAND2_X1 U268 ( .A1(n507), .A2(n506), .ZN(n253) );
  NAND2_X1 U270 ( .A1(\ML_int[2][16] ), .A2(n952), .ZN(n507) );
  NAND2_X1 U272 ( .A1(\ML_int[2][20] ), .A2(n967), .ZN(n506) );
  NAND2_X1 U273 ( .A1(n587), .A2(n586), .ZN(\ML_int[3][6] ) );
  NAND2_X1 U274 ( .A1(\ML_int[2][2] ), .A2(n952), .ZN(n587) );
  NAND2_X1 U275 ( .A1(\ML_int[2][6] ), .A2(n967), .ZN(n586) );
  NAND2_X1 U276 ( .A1(n321), .A2(n320), .ZN(n251) );
  NAND2_X1 U277 ( .A1(\ML_int[2][8] ), .A2(n953), .ZN(n321) );
  NAND2_X1 U278 ( .A1(\ML_int[2][12] ), .A2(n967), .ZN(n320) );
  NAND2_X1 U279 ( .A1(n521), .A2(net60893), .ZN(\ML_int[3][18] ) );
  NAND2_X1 U280 ( .A1(\ML_int[2][14] ), .A2(n953), .ZN(n521) );
  NAND2_X1 U282 ( .A1(\ML_int[2][18] ), .A2(n967), .ZN(net60893) );
  NAND2_X1 U283 ( .A1(n540), .A2(n539), .ZN(\ML_int[3][10] ) );
  NAND2_X1 U284 ( .A1(\ML_int[2][6] ), .A2(n953), .ZN(n540) );
  NAND2_X1 U285 ( .A1(\ML_int[2][10] ), .A2(n967), .ZN(n539) );
  NAND2_X1 U286 ( .A1(n538), .A2(n537), .ZN(\ML_int[3][11] ) );
  NAND2_X1 U287 ( .A1(\ML_int[2][7] ), .A2(n953), .ZN(n538) );
  NAND2_X1 U289 ( .A1(\ML_int[2][11] ), .A2(n967), .ZN(n537) );
  NAND2_X1 U290 ( .A1(n478), .A2(n479), .ZN(\MR_int[3][21] ) );
  NAND2_X1 U291 ( .A1(\MR_int[2][21] ), .A2(n954), .ZN(n478) );
  NAND2_X1 U292 ( .A1(\MR_int[2][25] ), .A2(n967), .ZN(n479) );
  NAND2_X1 U293 ( .A1(n556), .A2(n557), .ZN(\MR_int[3][9] ) );
  NAND2_X1 U295 ( .A1(\MR_int[2][9] ), .A2(n954), .ZN(n556) );
  NAND2_X1 U296 ( .A1(\MR_int[2][13] ), .A2(n967), .ZN(n557) );
  NAND2_X1 U297 ( .A1(n473), .A2(n474), .ZN(\ML_int[3][7] ) );
  NAND2_X1 U298 ( .A1(\ML_int[2][3] ), .A2(n955), .ZN(n474) );
  NAND2_X1 U300 ( .A1(\ML_int[2][7] ), .A2(n967), .ZN(n473) );
  NAND2_X1 U301 ( .A1(n141), .A2(n142), .ZN(\ML_int[3][15] ) );
  NAND2_X1 U302 ( .A1(\ML_int[2][11] ), .A2(n955), .ZN(n142) );
  NAND2_X1 U303 ( .A1(\ML_int[2][15] ), .A2(n967), .ZN(n141) );
  NAND2_X1 U304 ( .A1(n347), .A2(n346), .ZN(\MR_int[3][15] ) );
  NAND2_X1 U305 ( .A1(\MR_int[2][15] ), .A2(n955), .ZN(n346) );
  NAND2_X1 U306 ( .A1(\MR_int[2][19] ), .A2(n967), .ZN(n347) );
  NAND2_X1 U307 ( .A1(n300), .A2(n301), .ZN(\ML_int[3][5] ) );
  NAND2_X1 U308 ( .A1(\ML_int[2][1] ), .A2(n954), .ZN(n301) );
  NAND2_X1 U309 ( .A1(\ML_int[2][5] ), .A2(n967), .ZN(n300) );
  NAND2_X1 U310 ( .A1(n171), .A2(n1007), .ZN(n607) );
  NOR2_X1 U311 ( .A1(n968), .A2(n305), .ZN(n171) );
  AND2_X1 U312 ( .A1(n1018), .A2(n1044), .ZN(n205) );
  NAND2_X1 U313 ( .A1(\ML_int[3][25] ), .A2(n1008), .ZN(n488) );
  NAND2_X1 U314 ( .A1(n486), .A2(n487), .ZN(\ML_int[3][25] ) );
  NAND2_X1 U315 ( .A1(\ML_int[2][21] ), .A2(n951), .ZN(n487) );
  NAND2_X1 U316 ( .A1(\ML_int[2][25] ), .A2(n967), .ZN(n486) );
  NAND2_X1 U317 ( .A1(\ML_int[3][29] ), .A2(n1009), .ZN(n387) );
  NAND2_X1 U318 ( .A1(n390), .A2(n389), .ZN(\ML_int[3][29] ) );
  NAND2_X1 U319 ( .A1(\ML_int[2][25] ), .A2(n957), .ZN(n390) );
  NAND2_X1 U320 ( .A1(\ML_int[2][29] ), .A2(n967), .ZN(n389) );
  NAND2_X1 U321 ( .A1(n279), .A2(net60477), .ZN(\MR_int[3][22] ) );
  NAND2_X1 U322 ( .A1(n496), .A2(net61039), .ZN(\ML_int[3][17] ) );
  NAND2_X1 U323 ( .A1(n466), .A2(n465), .ZN(\ML_int[3][9] ) );
  NAND2_X1 U324 ( .A1(n348), .A2(n968), .ZN(n496) );
  NAND2_X1 U325 ( .A1(n410), .A2(n968), .ZN(n407) );
  INV_X1 U326 ( .A(n85), .ZN(n1042) );
  NAND2_X1 U327 ( .A1(\MR_int[3][13] ), .A2(n1007), .ZN(n127) );
  NAND2_X1 U328 ( .A1(\ML_int[2][24] ), .A2(n968), .ZN(n341) );
  NAND2_X1 U329 ( .A1(n250), .A2(n967), .ZN(n480) );
  AND2_X1 U330 ( .A1(\ML_int[2][0] ), .A2(n969), .ZN(\ML_int[3][0] ) );
  AND2_X1 U331 ( .A1(\ML_int[2][3] ), .A2(n967), .ZN(\ML_int[3][3] ) );
  AND2_X1 U332 ( .A1(\ML_int[2][1] ), .A2(n968), .ZN(\ML_int[3][1] ) );
  AND2_X1 U333 ( .A1(\ML_int[2][2] ), .A2(n969), .ZN(\ML_int[3][2] ) );
  OR2_X1 U334 ( .A1(n988), .A2(n1031), .ZN(n392) );
  AND2_X1 U335 ( .A1(\MR_int[3][29] ), .A2(n998), .ZN(\MR_int[4][29] ) );
  NOR2_X1 U336 ( .A1(n968), .A2(n305), .ZN(\MR_int[3][29] ) );
  AND2_X1 U338 ( .A1(n623), .A2(n624), .ZN(\MR_int[4][28] ) );
  NOR2_X1 U339 ( .A1(n1009), .A2(n968), .ZN(n624) );
  NAND2_X1 U340 ( .A1(\ML_int[2][5] ), .A2(n950), .ZN(n466) );
  BUF_X1 U341 ( .A(n173), .Z(n1010) );
  NAND2_X1 U342 ( .A1(n416), .A2(n415), .ZN(\ML_int[4][12] ) );
  NAND2_X1 U343 ( .A1(\ML_int[3][4] ), .A2(n993), .ZN(n416) );
  NAND2_X1 U344 ( .A1(n251), .A2(n1009), .ZN(n415) );
  NAND2_X1 U345 ( .A1(n395), .A2(n396), .ZN(\ML_int[4][13] ) );
  AND2_X1 U346 ( .A1(n355), .A2(n356), .ZN(n395) );
  NAND2_X1 U347 ( .A1(\ML_int[3][5] ), .A2(n994), .ZN(n396) );
  NAND2_X1 U348 ( .A1(n345), .A2(n357), .ZN(n355) );
  NAND2_X1 U349 ( .A1(n518), .A2(n519), .ZN(\ML_int[3][16] ) );
  NAND2_X1 U350 ( .A1(\ML_int[2][12] ), .A2(n956), .ZN(n519) );
  NAND2_X1 U351 ( .A1(\ML_int[2][16] ), .A2(n968), .ZN(n518) );
  NAND2_X1 U352 ( .A1(n220), .A2(n221), .ZN(n225) );
  AND2_X1 U353 ( .A1(n1015), .A2(n999), .ZN(n220) );
  NOR2_X1 U354 ( .A1(n392), .A2(n162), .ZN(n221) );
  NAND2_X1 U355 ( .A1(n958), .A2(net61436), .ZN(n162) );
  NAND2_X1 U356 ( .A1(n1014), .A2(n1044), .ZN(n676) );
  NAND2_X1 U357 ( .A1(n181), .A2(net61436), .ZN(n558) );
  NAND2_X1 U358 ( .A1(n332), .A2(n331), .ZN(n181) );
  NAND2_X1 U359 ( .A1(net61774), .A2(n1013), .ZN(n332) );
  NAND2_X1 U360 ( .A1(\MR_int[4][6] ), .A2(n1016), .ZN(n331) );
  NAND2_X1 U361 ( .A1(\MR_int[3][25] ), .A2(n1008), .ZN(n243) );
  INV_X1 U362 ( .A(\MR_int[2][30] ), .ZN(n1027) );
  NAND2_X1 U363 ( .A1(n552), .A2(n553), .ZN(\ML_int[3][14] ) );
  NAND2_X1 U366 ( .A1(\ML_int[2][10] ), .A2(n957), .ZN(n553) );
  NAND2_X1 U369 ( .A1(\ML_int[2][14] ), .A2(n969), .ZN(n552) );
  NAND2_X1 U371 ( .A1(n545), .A2(n546), .ZN(\MR_int[3][19] ) );
  NAND2_X1 U372 ( .A1(\MR_int[2][19] ), .A2(n956), .ZN(n546) );
  NAND2_X1 U373 ( .A1(\MR_int[2][23] ), .A2(n967), .ZN(n545) );
  NAND2_X1 U375 ( .A1(\MR_int[5][3] ), .A2(n549), .ZN(n576) );
  NAND2_X1 U376 ( .A1(n314), .A2(n315), .ZN(\MR_int[5][3] ) );
  NAND2_X1 U377 ( .A1(\MR_int[4][3] ), .A2(n1016), .ZN(n314) );
  NAND2_X1 U378 ( .A1(\MR_int[4][19] ), .A2(n1013), .ZN(n315) );
  NAND2_X1 U379 ( .A1(n272), .A2(n273), .ZN(n499) );
  NAND2_X1 U380 ( .A1(n1024), .A2(n412), .ZN(n272) );
  INV_X1 U381 ( .A(n690), .ZN(n1024) );
  NAND2_X1 U382 ( .A1(\MR_int[4][25] ), .A2(n1013), .ZN(n412) );
  BUF_X1 U383 ( .A(\temp_int_SH[4] ), .Z(n1018) );
  AND2_X1 U384 ( .A1(\MR_int[3][25] ), .A2(n999), .ZN(\MR_int[4][25] ) );
  NAND2_X1 U385 ( .A1(\ML_int[7][0] ), .A2(n947), .ZN(n502) );
  NOR2_X1 U386 ( .A1(n325), .A2(n88), .ZN(\ML_int[7][0] ) );
  NAND2_X1 U387 ( .A1(n235), .A2(n622), .ZN(n447) );
  AND2_X1 U388 ( .A1(\ML_int[4][12] ), .A2(n948), .ZN(n235) );
  NAND2_X1 U390 ( .A1(\ML_int[2][20] ), .A2(n950), .ZN(n342) );
  NAND2_X1 U391 ( .A1(\ML_int[2][23] ), .A2(n950), .ZN(n481) );
  NAND2_X1 U392 ( .A1(\MR_int[3][5] ), .A2(n991), .ZN(n128) );
  NAND2_X1 U393 ( .A1(\ML_int[7][2] ), .A2(n946), .ZN(n577) );
  NOR2_X1 U394 ( .A1(n325), .A2(n86), .ZN(\ML_int[7][2] ) );
  NAND2_X1 U395 ( .A1(\ML_int[7][4] ), .A2(n946), .ZN(n340) );
  NOR2_X1 U396 ( .A1(n325), .A2(n83), .ZN(\ML_int[7][4] ) );
  NAND2_X1 U397 ( .A1(net141573), .A2(n1008), .ZN(n83) );
  NAND2_X1 U398 ( .A1(\ML_int[7][5] ), .A2(n946), .ZN(n559) );
  NOR2_X1 U399 ( .A1(n82), .A2(n325), .ZN(\ML_int[7][5] ) );
  NAND2_X1 U400 ( .A1(\ML_int[7][6] ), .A2(n946), .ZN(n461) );
  NOR2_X1 U401 ( .A1(n325), .A2(n81), .ZN(\ML_int[7][6] ) );
  NAND2_X1 U402 ( .A1(\ML_int[7][10] ), .A2(n946), .ZN(n585) );
  AND2_X1 U403 ( .A1(\ML_int[4][10] ), .A2(n622), .ZN(\ML_int[7][10] ) );
  NAND2_X1 U404 ( .A1(\ML_int[7][14] ), .A2(n946), .ZN(n569) );
  AND2_X1 U405 ( .A1(\ML_int[4][14] ), .A2(n622), .ZN(\ML_int[7][14] ) );
  NAND2_X1 U406 ( .A1(\ML_int[7][1] ), .A2(n947), .ZN(n611) );
  NOR2_X1 U407 ( .A1(n325), .A2(n87), .ZN(\ML_int[7][1] ) );
  NAND2_X1 U408 ( .A1(n725), .A2(n1013), .ZN(n448) );
  NAND2_X1 U409 ( .A1(n522), .A2(n523), .ZN(\MR_int[4][20] ) );
  NAND2_X1 U410 ( .A1(n384), .A2(n622), .ZN(n455) );
  AND2_X1 U411 ( .A1(\ML_int[4][15] ), .A2(n948), .ZN(n384) );
  NAND2_X1 U412 ( .A1(\ML_int[2][24] ), .A2(n951), .ZN(n418) );
  NAND2_X1 U413 ( .A1(\MR_int[2][8] ), .A2(n951), .ZN(n406) );
  NAND2_X1 U414 ( .A1(\ML_int[3][21] ), .A2(n992), .ZN(n386) );
  NAND2_X1 U415 ( .A1(\ML_int[7][28] ), .A2(n946), .ZN(n318) );
  NAND2_X1 U416 ( .A1(n375), .A2(n376), .ZN(\ML_int[7][28] ) );
  NAND2_X1 U417 ( .A1(\ML_int[4][12] ), .A2(n377), .ZN(n375) );
  NAND2_X1 U418 ( .A1(\ML_int[4][28] ), .A2(n252), .ZN(n376) );
  NAND2_X1 U419 ( .A1(n738), .A2(n739), .ZN(n454) );
  NAND2_X1 U420 ( .A1(n627), .A2(n628), .ZN(n738) );
  NOR2_X1 U421 ( .A1(n1014), .A2(net61266), .ZN(n739) );
  NAND2_X1 U422 ( .A1(\MR_int[3][16] ), .A2(n992), .ZN(n627) );
  NAND2_X1 U423 ( .A1(\MR_int[4][22] ), .A2(n189), .ZN(n428) );
  NOR2_X1 U424 ( .A1(n1014), .A2(net61266), .ZN(n189) );
  BUF_X1 U425 ( .A(n173), .Z(n1011) );
  NAND2_X1 U426 ( .A1(n337), .A2(n338), .ZN(\MR_int[4][13] ) );
  NAND2_X1 U427 ( .A1(net141562), .A2(n991), .ZN(n337) );
  NAND2_X1 U428 ( .A1(\MR_int[3][21] ), .A2(n1008), .ZN(n338) );
  NAND2_X1 U429 ( .A1(n800), .A2(n801), .ZN(n451) );
  NAND2_X1 U430 ( .A1(n574), .A2(n575), .ZN(n801) );
  NOR2_X1 U431 ( .A1(net60660), .A2(n1013), .ZN(n800) );
  NAND2_X1 U432 ( .A1(\MR_int[3][26] ), .A2(n1008), .ZN(n574) );
  NAND2_X1 U433 ( .A1(n200), .A2(n505), .ZN(\ML_int[2][9] ) );
  NAND2_X1 U434 ( .A1(\MR_int[4][8] ), .A2(n257), .ZN(n255) );
  AND2_X1 U435 ( .A1(n1018), .A2(n237), .ZN(n257) );
  NAND2_X1 U436 ( .A1(n406), .A2(n407), .ZN(\MR_int[3][8] ) );
  NAND2_X1 U437 ( .A1(\MR_int[4][4] ), .A2(n214), .ZN(n212) );
  AND2_X1 U438 ( .A1(n1018), .A2(n273), .ZN(n214) );
  NAND2_X1 U439 ( .A1(net60588), .A2(net60589), .ZN(\MR_int[3][14] ) );
  NAND2_X1 U440 ( .A1(n660), .A2(n575), .ZN(\MR_int[4][18] ) );
  NAND2_X1 U441 ( .A1(\MR_int[3][26] ), .A2(n1008), .ZN(n660) );
  NAND2_X1 U442 ( .A1(n605), .A2(n604), .ZN(\MR_int[4][19] ) );
  NAND2_X1 U443 ( .A1(\MR_int[3][27] ), .A2(n1008), .ZN(n605) );
  NAND2_X1 U444 ( .A1(n156), .A2(n157), .ZN(n572) );
  NAND2_X1 U445 ( .A1(n522), .A2(n523), .ZN(n156) );
  NOR2_X1 U446 ( .A1(n1013), .A2(net60660), .ZN(n157) );
  NAND2_X1 U447 ( .A1(\ML_int[5][26] ), .A2(n493), .ZN(n525) );
  NAND2_X1 U449 ( .A1(n299), .A2(n298), .ZN(\ML_int[5][26] ) );
  NAND2_X1 U450 ( .A1(\ML_int[4][10] ), .A2(n1017), .ZN(n299) );
  NAND2_X1 U451 ( .A1(\ML_int[4][26] ), .A2(n1012), .ZN(n298) );
  NAND2_X1 U452 ( .A1(n279), .A2(net60477), .ZN(n727) );
  NAND2_X1 U453 ( .A1(n547), .A2(n548), .ZN(\MR_int[2][17] ) );
  NAND2_X1 U454 ( .A1(net61755), .A2(n349), .ZN(\MR_int[4][6] ) );
  NAND2_X1 U455 ( .A1(\MR_int[3][6] ), .A2(n991), .ZN(n349) );
  NAND2_X1 U456 ( .A1(\MR_int[3][14] ), .A2(n1007), .ZN(net61755) );
  AND2_X1 U457 ( .A1(n1017), .A2(n85), .ZN(n377) );
  AND2_X1 U458 ( .A1(n1017), .A2(n85), .ZN(n736) );
  NAND2_X1 U459 ( .A1(n163), .A2(n164), .ZN(n568) );
  NAND2_X1 U460 ( .A1(n225), .A2(n760), .ZN(n164) );
  NAND2_X1 U461 ( .A1(n1017), .A2(n306), .ZN(n760) );
  NAND2_X1 U462 ( .A1(\MR_int[4][14] ), .A2(n170), .ZN(n667) );
  AND2_X1 U463 ( .A1(n1017), .A2(net61436), .ZN(n170) );
  NAND2_X1 U464 ( .A1(net60588), .A2(net60589), .ZN(n669) );
  NAND2_X1 U465 ( .A1(\ML_int[5][21] ), .A2(net61624), .ZN(n427) );
  NAND2_X1 U466 ( .A1(n124), .A2(n125), .ZN(\ML_int[5][21] ) );
  AND2_X1 U467 ( .A1(n85), .A2(n948), .ZN(net61624) );
  NAND2_X1 U468 ( .A1(\ML_int[4][21] ), .A2(n1012), .ZN(n124) );
  NAND2_X1 U469 ( .A1(\ML_int[5][30] ), .A2(n421), .ZN(n529) );
  NAND2_X1 U470 ( .A1(n714), .A2(n715), .ZN(\ML_int[5][30] ) );
  AND2_X1 U471 ( .A1(n85), .A2(n948), .ZN(n421) );
  NAND2_X1 U472 ( .A1(\ML_int[4][30] ), .A2(n1012), .ZN(n714) );
  NAND2_X1 U473 ( .A1(\MR_int[4][12] ), .A2(n241), .ZN(n723) );
  AND2_X1 U474 ( .A1(n1017), .A2(n405), .ZN(n241) );
  NAND2_X1 U475 ( .A1(n554), .A2(n555), .ZN(\MR_int[3][11] ) );
  NAND2_X1 U476 ( .A1(\MR_int[2][11] ), .A2(n957), .ZN(n554) );
  NAND2_X1 U477 ( .A1(\MR_int[2][15] ), .A2(n968), .ZN(n555) );
  NAND2_X1 U478 ( .A1(n558), .A2(n559), .ZN(B[5]) );
  NAND2_X1 U479 ( .A1(n460), .A2(n461), .ZN(B[6]) );
  NAND2_X1 U480 ( .A1(n178), .A2(n255), .ZN(B[7]) );
  AND2_X1 U481 ( .A1(\ML_int[5][31] ), .A2(n378), .ZN(B[31]) );
  NAND2_X1 U482 ( .A1(n584), .A2(n585), .ZN(B[10]) );
  NAND2_X1 U483 ( .A1(n514), .A2(n515), .ZN(B[23]) );
  NAND2_X1 U484 ( .A1(n667), .A2(n668), .ZN(B[13]) );
  NAND2_X1 U485 ( .A1(n446), .A2(n447), .ZN(B[12]) );
  NAND2_X1 U486 ( .A1(n455), .A2(n454), .ZN(B[15]) );
  NAND2_X1 U487 ( .A1(n450), .A2(n451), .ZN(B[17]) );
  NAND2_X1 U488 ( .A1(n336), .A2(n335), .ZN(B[25]) );
  NAND2_X1 U489 ( .A1(n525), .A2(n524), .ZN(B[26]) );
  OR2_X1 U490 ( .A1(n271), .A2(n948), .ZN(n335) );
  NAND2_X1 U491 ( .A1(n1044), .A2(n274), .ZN(n271) );
  NOR2_X1 U492 ( .A1(n1014), .A2(n385), .ZN(n274) );
  NAND2_X1 U494 ( .A1(n998), .A2(\MR_int[3][26] ), .ZN(n385) );
  OR2_X1 U495 ( .A1(n358), .A2(n359), .ZN(n435) );
  NAND2_X1 U496 ( .A1(n223), .A2(n1016), .ZN(n358) );
  NAND2_X1 U497 ( .A1(net61842), .A2(n604), .ZN(n223) );
  NAND2_X1 U498 ( .A1(n236), .A2(n1008), .ZN(net61842) );
  OR2_X1 U499 ( .A1(n388), .A2(net60660), .ZN(n524) );
  OR2_X1 U500 ( .A1(n197), .A2(n1015), .ZN(n388) );
  NAND2_X1 U501 ( .A1(n726), .A2(n995), .ZN(n197) );
  OR2_X1 U502 ( .A1(n324), .A2(n359), .ZN(n401) );
  OR2_X1 U503 ( .A1(n1026), .A2(n1014), .ZN(n324) );
  INV_X1 U504 ( .A(\MR_int[4][28] ), .ZN(n1026) );
  OR2_X1 U505 ( .A1(n207), .A2(n208), .ZN(n319) );
  OR2_X1 U506 ( .A1(n1025), .A2(n1014), .ZN(n207) );
  INV_X1 U507 ( .A(\MR_int[4][29] ), .ZN(n1025) );
  NAND2_X1 U508 ( .A1(\ML_int[7][9] ), .A2(n946), .ZN(n594) );
  AND2_X1 U509 ( .A1(\ML_int[4][9] ), .A2(n622), .ZN(\ML_int[7][9] ) );
  AND2_X1 U510 ( .A1(net60718), .A2(n168), .ZN(n668) );
  OR2_X1 U511 ( .A1(n476), .A2(n180), .ZN(n168) );
  NAND2_X1 U512 ( .A1(\ML_int[7][13] ), .A2(n946), .ZN(net60718) );
  NAND2_X1 U513 ( .A1(\MR_int[4][30] ), .A2(n1012), .ZN(n180) );
  OR2_X1 U514 ( .A1(n1017), .A2(n476), .ZN(n737) );
  AND2_X1 U515 ( .A1(n724), .A2(n532), .ZN(n666) );
  NAND2_X1 U516 ( .A1(\ML_int[4][11] ), .A2(n211), .ZN(n532) );
  OR2_X1 U517 ( .A1(n208), .A2(n592), .ZN(n724) );
  AND2_X1 U518 ( .A1(n622), .A2(n948), .ZN(n211) );
  NAND2_X1 U519 ( .A1(n308), .A2(n307), .ZN(\MR_int[3][12] ) );
  NAND2_X1 U520 ( .A1(n410), .A2(n958), .ZN(n307) );
  NAND2_X1 U521 ( .A1(\MR_int[2][16] ), .A2(n969), .ZN(n308) );
  BUF_X1 U522 ( .A(n965), .Z(n963) );
  BUF_X1 U523 ( .A(n965), .Z(n964) );
  BUF_X1 U524 ( .A(n966), .Z(n962) );
  BUF_X1 U525 ( .A(n966), .Z(n961) );
  BUF_X1 U526 ( .A(n1005), .Z(n1004) );
  BUF_X1 U527 ( .A(n1005), .Z(n1003) );
  BUF_X1 U528 ( .A(n1006), .Z(n1001) );
  BUF_X1 U529 ( .A(n1006), .Z(n1002) );
  NAND2_X1 U530 ( .A1(net61331), .A2(n439), .ZN(\MR_int[3][10] ) );
  NAND2_X1 U531 ( .A1(\MR_int[2][10] ), .A2(n958), .ZN(n439) );
  NAND2_X1 U532 ( .A1(\MR_int[2][14] ), .A2(n967), .ZN(net61331) );
  NAND2_X1 U533 ( .A1(n1020), .A2(n401), .ZN(B[27]) );
  NAND2_X1 U534 ( .A1(n723), .A2(n666), .ZN(B[11]) );
  NAND2_X1 U535 ( .A1(n427), .A2(n428), .ZN(B[21]) );
  AND2_X1 U536 ( .A1(n583), .A2(n213), .ZN(n696) );
  NAND2_X1 U537 ( .A1(\MR_int[4][20] ), .A2(n201), .ZN(n213) );
  NAND2_X1 U538 ( .A1(\ML_int[7][3] ), .A2(n946), .ZN(n583) );
  AND2_X1 U539 ( .A1(n1015), .A2(n549), .ZN(n201) );
  AND2_X1 U540 ( .A1(n477), .A2(n256), .ZN(n178) );
  OR2_X1 U541 ( .A1(n359), .A2(n449), .ZN(n256) );
  NAND2_X1 U542 ( .A1(\ML_int[7][7] ), .A2(n946), .ZN(n477) );
  NAND2_X1 U543 ( .A1(n730), .A2(n175), .ZN(n449) );
  AND2_X1 U544 ( .A1(n708), .A2(n709), .ZN(n446) );
  NAND2_X1 U545 ( .A1(\MR_int[4][13] ), .A2(n204), .ZN(n708) );
  OR2_X1 U546 ( .A1(n359), .A2(n456), .ZN(n709) );
  AND2_X1 U547 ( .A1(n1018), .A2(n237), .ZN(n204) );
  AND2_X1 U548 ( .A1(n578), .A2(n579), .ZN(n224) );
  NAND2_X1 U549 ( .A1(\MR_int[3][17] ), .A2(n997), .ZN(n579) );
  NAND2_X1 U550 ( .A1(\MR_int[3][25] ), .A2(n1008), .ZN(n578) );
  NAND2_X1 U551 ( .A1(n1019), .A2(n611), .ZN(B[1]) );
  NAND2_X1 U552 ( .A1(n318), .A2(n319), .ZN(B[28]) );
  AND2_X1 U553 ( .A1(n85), .A2(n948), .ZN(n378) );
  NAND2_X1 U554 ( .A1(n131), .A2(n132), .ZN(\ML_int[5][31] ) );
  NAND2_X1 U555 ( .A1(\ML_int[4][31] ), .A2(n1012), .ZN(n131) );
  NAND2_X1 U556 ( .A1(\ML_int[4][15] ), .A2(n1016), .ZN(n132) );
  INV_X1 U559 ( .A(n295), .ZN(n1022) );
  OAI21_X1 U560 ( .B1(n1014), .B2(n673), .A(n744), .ZN(n295) );
  NAND2_X1 U561 ( .A1(\MR_int[3][9] ), .A2(n745), .ZN(n744) );
  NAND2_X1 U562 ( .A1(\MR_int[3][1] ), .A2(n996), .ZN(n673) );
  OR2_X1 U563 ( .A1(n802), .A2(n803), .ZN(n233) );
  NAND2_X1 U564 ( .A1(n237), .A2(n1013), .ZN(n803) );
  NAND2_X1 U566 ( .A1(\MR_int[3][26] ), .A2(n992), .ZN(n802) );
  NAND2_X1 U567 ( .A1(\MR_int[4][10] ), .A2(n234), .ZN(n232) );
  AND2_X1 U568 ( .A1(n1017), .A2(n261), .ZN(n234) );
  INV_X1 U569 ( .A(n459), .ZN(n1041) );
  INV_X1 U570 ( .A(n691), .ZN(n1019) );
  AOI21_X1 U571 ( .B1(n589), .B2(n588), .A(n476), .ZN(n691) );
  NAND2_X1 U572 ( .A1(\MR_int[4][18] ), .A2(n1013), .ZN(n589) );
  NAND2_X1 U573 ( .A1(\MR_int[4][2] ), .A2(n1016), .ZN(n588) );
  AND2_X1 U574 ( .A1(\SHMAG[5] ), .A2(n948), .ZN(n85) );
  NAND2_X1 U575 ( .A1(n106), .A2(n947), .ZN(net61465) );
  NAND4_X1 U576 ( .A1(n109), .A2(n110), .A3(n107), .A4(n108), .ZN(n106) );
  NAND2_X1 U577 ( .A1(net61465), .A2(net141444), .ZN(net135734) );
  NOR2_X1 U578 ( .A1(\SHMAG[5] ), .A2(n947), .ZN(net61436) );
  NAND2_X1 U579 ( .A1(n89), .A2(n96), .ZN(\temp_int_SH[0] ) );
  BUF_X1 U580 ( .A(n1046), .Z(n946) );
  BUF_X1 U581 ( .A(n1046), .Z(n947) );
  BUF_X1 U583 ( .A(n1046), .Z(n948) );
  NOR2_X1 U584 ( .A1(n947), .A2(\SHMAG[5] ), .ZN(n237) );
  OAI221_X1 U585 ( .B1(n1022), .B2(n476), .C1(n224), .C2(n737), .A(n502), .ZN(
        B[0]) );
  NOR2_X1 U586 ( .A1(n947), .A2(\SHMAG[5] ), .ZN(n549) );
  NOR2_X1 U587 ( .A1(n947), .A2(\SHMAG[5] ), .ZN(n273) );
  NOR2_X1 U588 ( .A1(n947), .A2(\SHMAG[5] ), .ZN(n261) );
  NAND2_X1 U589 ( .A1(net61465), .A2(net141444), .ZN(net61851) );
  NAND4_X1 U590 ( .A1(n285), .A2(n286), .A3(n284), .A4(n270), .ZN(net60578) );
  AND2_X1 U591 ( .A1(net60450), .A2(n104), .ZN(n286) );
  NOR2_X1 U592 ( .A1(net60750), .A2(net60751), .ZN(n285) );
  NOR2_X1 U593 ( .A1(net61363), .A2(net61364), .ZN(n284) );
  INV_X1 U594 ( .A(\SHMAG[5] ), .ZN(n1044) );
  NOR2_X1 U595 ( .A1(\SHMAG[5] ), .A2(n947), .ZN(n306) );
  NAND2_X1 U596 ( .A1(net61465), .A2(net141444), .ZN(n729) );
  NOR2_X1 U597 ( .A1(n947), .A2(\SHMAG[5] ), .ZN(n405) );
  NOR2_X1 U598 ( .A1(n1014), .A2(\SHMAG[5] ), .ZN(n391) );
  NOR2_X1 U599 ( .A1(net65464), .A2(net65465), .ZN(n270) );
  NOR2_X1 U600 ( .A1(net61363), .A2(net61364), .ZN(n100) );
  NAND2_X1 U602 ( .A1(n656), .A2(n947), .ZN(n89) );
  NAND4_X1 U603 ( .A1(n109), .A2(n110), .A3(n107), .A4(n108), .ZN(n656) );
  AND2_X1 U604 ( .A1(n96), .A2(n89), .ZN(net141501) );
  NAND2_X1 U605 ( .A1(net61465), .A2(n90), .ZN(\temp_int_SH[4] ) );
  NOR2_X1 U606 ( .A1(net65464), .A2(net65465), .ZN(n98) );
  OR2_X1 U607 ( .A1(\SHMAG[5] ), .A2(n948), .ZN(n476) );
  NAND2_X1 U609 ( .A1(n228), .A2(n1009), .ZN(n523) );
  NOR2_X1 U610 ( .A1(n968), .A2(n215), .ZN(n228) );
  AND2_X1 U611 ( .A1(n570), .A2(n571), .ZN(n215) );
  NAND2_X1 U612 ( .A1(\MR_int[2][26] ), .A2(n968), .ZN(net60477) );
  NAND2_X1 U613 ( .A1(\MR_int[1][19] ), .A2(n988), .ZN(n548) );
  NAND2_X1 U614 ( .A1(\MR_int[2][18] ), .A2(n969), .ZN(net60588) );
  NAND2_X1 U615 ( .A1(n712), .A2(n713), .ZN(\MR_int[2][27] ) );
  NAND2_X1 U616 ( .A1(\MR_int[1][27] ), .A2(n971), .ZN(n713) );
  NAND2_X1 U617 ( .A1(\ML_int[1][30] ), .A2(n986), .ZN(n712) );
  NAND2_X1 U618 ( .A1(n147), .A2(n148), .ZN(\MR_int[3][25] ) );
  NAND2_X1 U619 ( .A1(\MR_int[2][25] ), .A2(n952), .ZN(n148) );
  NAND2_X1 U620 ( .A1(\MR_int[2][29] ), .A2(n967), .ZN(n147) );
  NAND2_X1 U622 ( .A1(n597), .A2(n598), .ZN(\MR_int[2][29] ) );
  NAND2_X1 U623 ( .A1(\ML_int[1][9] ), .A2(n987), .ZN(n200) );
  NAND2_X1 U624 ( .A1(\ML_int[1][17] ), .A2(n988), .ZN(n457) );
  NOR2_X1 U625 ( .A1(\SHMAG[5] ), .A2(n15), .ZN(\MR_int[7][29] ) );
  OR2_X1 U626 ( .A1(n1014), .A2(n743), .ZN(n15) );
  NAND2_X1 U627 ( .A1(n997), .A2(n155), .ZN(n743) );
  OR2_X1 U628 ( .A1(n948), .A2(\SHMAG[5] ), .ZN(net60660) );
  NAND2_X1 U629 ( .A1(\MR_int[1][31] ), .A2(n986), .ZN(n598) );
  NAND2_X1 U630 ( .A1(\MR_int[1][30] ), .A2(n987), .ZN(n570) );
  NAND2_X1 U631 ( .A1(\ML_int[1][19] ), .A2(n988), .ZN(n352) );
  NAND2_X1 U632 ( .A1(\ML_int[1][7] ), .A2(n970), .ZN(n505) );
  OR2_X1 U633 ( .A1(n948), .A2(\SHMAG[5] ), .ZN(n359) );
  NAND2_X1 U634 ( .A1(n264), .A2(n949), .ZN(net61039) );
  NAND2_X1 U635 ( .A1(n344), .A2(n343), .ZN(\ML_int[2][15] ) );
  NAND2_X1 U636 ( .A1(n728), .A2(n971), .ZN(n344) );
  NAND2_X1 U637 ( .A1(n988), .A2(\MR_int[1][14] ), .ZN(n343) );
  NAND2_X1 U638 ( .A1(\ML_int[1][19] ), .A2(n970), .ZN(n459) );
  NAND2_X1 U639 ( .A1(\MR_int[1][17] ), .A2(n970), .ZN(n547) );
  NAND2_X1 U640 ( .A1(n457), .A2(n302), .ZN(n348) );
  NAND2_X1 U641 ( .A1(n492), .A2(n334), .ZN(\ML_int[2][8] ) );
  NAND2_X1 U642 ( .A1(\ML_int[1][6] ), .A2(n971), .ZN(n492) );
  NAND2_X1 U643 ( .A1(\MR_int[2][22] ), .A2(n949), .ZN(n279) );
  NAND2_X1 U644 ( .A1(n608), .A2(n609), .ZN(\MR_int[2][21] ) );
  NAND2_X1 U645 ( .A1(\MR_int[1][21] ), .A2(n974), .ZN(n608) );
  NAND2_X1 U646 ( .A1(n601), .A2(n987), .ZN(n609) );
  NAND2_X1 U647 ( .A1(net61783), .A2(net61782), .ZN(\ML_int[2][20] ) );
  NAND2_X1 U648 ( .A1(\ML_int[1][18] ), .A2(n975), .ZN(net61783) );
  NAND2_X1 U649 ( .A1(\ML_int[1][20] ), .A2(n987), .ZN(net61782) );
  NAND2_X1 U650 ( .A1(n404), .A2(n403), .ZN(\ML_int[2][16] ) );
  NAND2_X1 U651 ( .A1(\ML_int[1][14] ), .A2(n975), .ZN(n404) );
  NAND2_X1 U652 ( .A1(\ML_int[1][16] ), .A2(n987), .ZN(n403) );
  NAND2_X1 U653 ( .A1(n599), .A2(n600), .ZN(\MR_int[2][24] ) );
  NAND2_X1 U654 ( .A1(\MR_int[1][24] ), .A2(n975), .ZN(n599) );
  NAND2_X1 U655 ( .A1(\MR_int[1][26] ), .A2(n987), .ZN(n600) );
  NAND2_X1 U656 ( .A1(n595), .A2(n596), .ZN(\MR_int[2][19] ) );
  NAND2_X1 U657 ( .A1(\MR_int[1][19] ), .A2(n974), .ZN(n595) );
  NAND2_X1 U658 ( .A1(\MR_int[1][21] ), .A2(n987), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n351), .A2(n350), .ZN(\ML_int[2][11] ) );
  NAND2_X1 U660 ( .A1(\ML_int[1][9] ), .A2(n976), .ZN(n351) );
  NAND2_X1 U661 ( .A1(\ML_int[1][11] ), .A2(n987), .ZN(n350) );
  NAND2_X1 U662 ( .A1(n543), .A2(n544), .ZN(\MR_int[2][25] ) );
  NAND2_X1 U663 ( .A1(\MR_int[1][25] ), .A2(n975), .ZN(n543) );
  NAND2_X1 U664 ( .A1(\MR_int[1][27] ), .A2(n987), .ZN(n544) );
  NAND2_X1 U665 ( .A1(n398), .A2(n397), .ZN(\ML_int[2][10] ) );
  NAND2_X1 U666 ( .A1(\MR_int[1][7] ), .A2(n976), .ZN(n398) );
  NAND2_X1 U667 ( .A1(\ML_int[1][10] ), .A2(n987), .ZN(n397) );
  NAND2_X1 U668 ( .A1(n542), .A2(net60763), .ZN(\MR_int[2][16] ) );
  NAND2_X1 U669 ( .A1(\MR_int[1][16] ), .A2(n976), .ZN(n542) );
  NAND2_X1 U670 ( .A1(\MR_int[1][18] ), .A2(n987), .ZN(net60763) );
  NAND2_X1 U671 ( .A1(n121), .A2(n122), .ZN(\ML_int[2][23] ) );
  NAND2_X1 U672 ( .A1(\ML_int[1][21] ), .A2(n972), .ZN(n122) );
  NAND2_X1 U673 ( .A1(\ML_int[1][23] ), .A2(n986), .ZN(n121) );
  NAND2_X1 U674 ( .A1(n283), .A2(n282), .ZN(\MR_int[2][14] ) );
  NAND2_X1 U675 ( .A1(\MR_int[1][14] ), .A2(n972), .ZN(n282) );
  NAND2_X1 U676 ( .A1(\MR_int[1][16] ), .A2(n987), .ZN(n283) );
  NAND2_X1 U677 ( .A1(n581), .A2(net60604), .ZN(\MR_int[2][15] ) );
  NAND2_X1 U678 ( .A1(\ML_int[1][16] ), .A2(n973), .ZN(net60604) );
  NAND2_X1 U679 ( .A1(\MR_int[1][17] ), .A2(n986), .ZN(n581) );
  NAND2_X1 U680 ( .A1(n482), .A2(n483), .ZN(\ML_int[2][12] ) );
  NAND2_X1 U681 ( .A1(\ML_int[1][10] ), .A2(n973), .ZN(n483) );
  NAND2_X1 U682 ( .A1(\ML_int[1][12] ), .A2(n987), .ZN(n482) );
  NAND2_X1 U683 ( .A1(n706), .A2(n707), .ZN(\MR_int[2][23] ) );
  NAND2_X1 U684 ( .A1(n601), .A2(n972), .ZN(n707) );
  NAND2_X1 U685 ( .A1(\MR_int[1][25] ), .A2(n987), .ZN(n706) );
  NAND2_X1 U686 ( .A1(n508), .A2(n509), .ZN(\ML_int[2][14] ) );
  NAND2_X1 U687 ( .A1(\ML_int[1][12] ), .A2(n973), .ZN(n509) );
  NAND2_X1 U688 ( .A1(\ML_int[1][14] ), .A2(n988), .ZN(n508) );
  NAND2_X1 U689 ( .A1(n452), .A2(n453), .ZN(\ML_int[2][25] ) );
  NAND2_X1 U690 ( .A1(\ML_int[1][23] ), .A2(n974), .ZN(n453) );
  NAND2_X1 U691 ( .A1(\ML_int[1][25] ), .A2(n987), .ZN(n452) );
  NAND2_X1 U692 ( .A1(n440), .A2(n441), .ZN(\ML_int[2][7] ) );
  NAND2_X1 U693 ( .A1(\ML_int[1][5] ), .A2(n974), .ZN(n441) );
  NAND2_X1 U694 ( .A1(\ML_int[1][7] ), .A2(n987), .ZN(n440) );
  NAND2_X1 U695 ( .A1(n393), .A2(n394), .ZN(\ML_int[2][6] ) );
  NAND2_X1 U696 ( .A1(\MR_int[1][3] ), .A2(n973), .ZN(n394) );
  NAND2_X1 U697 ( .A1(\ML_int[1][6] ), .A2(n986), .ZN(n393) );
  NAND2_X1 U698 ( .A1(n699), .A2(n700), .ZN(\ML_int[2][5] ) );
  NAND2_X1 U699 ( .A1(\ML_int[1][3] ), .A2(n972), .ZN(n700) );
  NAND2_X1 U700 ( .A1(\ML_int[1][5] ), .A2(n987), .ZN(n699) );
  OR2_X1 U701 ( .A1(n948), .A2(\SHMAG[5] ), .ZN(net61266) );
  NAND2_X1 U702 ( .A1(n153), .A2(n154), .ZN(\MR_int[2][2] ) );
  NAND2_X1 U703 ( .A1(\MR_int[1][2] ), .A2(n977), .ZN(n154) );
  AND2_X1 U704 ( .A1(n598), .A2(n597), .ZN(n305) );
  NAND2_X1 U705 ( .A1(n530), .A2(net60869), .ZN(\ML_int[2][4] ) );
  NAND2_X1 U706 ( .A1(\ML_int[1][2] ), .A2(n976), .ZN(n530) );
  NAND2_X1 U707 ( .A1(\ML_int[1][4] ), .A2(n986), .ZN(net60869) );
  NAND2_X1 U708 ( .A1(n517), .A2(n516), .ZN(\ML_int[3][13] ) );
  NAND2_X1 U709 ( .A1(\ML_int[2][9] ), .A2(n951), .ZN(n517) );
  NAND2_X1 U710 ( .A1(\ML_int[2][13] ), .A2(n968), .ZN(n516) );
  NAND2_X1 U711 ( .A1(\MR_int[1][4] ), .A2(n986), .ZN(n153) );
  NAND2_X1 U712 ( .A1(\ML_int[1][17] ), .A2(n970), .ZN(n353) );
  NAND2_X1 U713 ( .A1(n571), .A2(n570), .ZN(n623) );
  NAND2_X1 U714 ( .A1(n195), .A2(n196), .ZN(\ML_int[2][2] ) );
  NAND2_X1 U715 ( .A1(\ML_int[1][0] ), .A2(n977), .ZN(n196) );
  NAND2_X1 U716 ( .A1(\ML_int[1][2] ), .A2(n986), .ZN(n195) );
  NAND2_X1 U717 ( .A1(n511), .A2(n510), .ZN(\ML_int[3][21] ) );
  NAND2_X1 U718 ( .A1(\ML_int[2][17] ), .A2(n954), .ZN(n511) );
  AOI22_X1 U719 ( .A1(n731), .A2(\ML_int[1][21] ), .B1(n1041), .B2(n968), .ZN(
        n510) );
  NAND2_X1 U720 ( .A1(n457), .A2(n302), .ZN(\ML_int[2][17] ) );
  NAND2_X1 U721 ( .A1(n333), .A2(n334), .ZN(\MR_int[2][5] ) );
  NAND2_X1 U722 ( .A1(\MR_int[1][5] ), .A2(n977), .ZN(n333) );
  NAND2_X1 U723 ( .A1(n566), .A2(n567), .ZN(\MR_int[3][20] ) );
  NAND2_X1 U724 ( .A1(\MR_int[2][20] ), .A2(n955), .ZN(n566) );
  NAND2_X1 U725 ( .A1(\MR_int[2][24] ), .A2(n967), .ZN(n567) );
  NAND2_X1 U726 ( .A1(n535), .A2(n536), .ZN(\MR_int[3][18] ) );
  NAND2_X1 U727 ( .A1(net61353), .A2(n956), .ZN(n535) );
  NAND2_X1 U728 ( .A1(\MR_int[2][22] ), .A2(n967), .ZN(n536) );
  NAND2_X1 U729 ( .A1(n497), .A2(n498), .ZN(\MR_int[2][8] ) );
  NAND2_X1 U730 ( .A1(\MR_int[1][8] ), .A2(n978), .ZN(n497) );
  NAND2_X1 U731 ( .A1(\MR_int[1][10] ), .A2(n986), .ZN(n498) );
  NAND2_X1 U733 ( .A1(n326), .A2(n327), .ZN(\ML_int[2][18] ) );
  NAND2_X1 U735 ( .A1(\MR_int[1][15] ), .A2(n977), .ZN(n327) );
  NAND2_X1 U736 ( .A1(\ML_int[1][18] ), .A2(n986), .ZN(n326) );
  NAND2_X1 U737 ( .A1(n591), .A2(n590), .ZN(\MR_int[3][16] ) );
  NAND2_X1 U738 ( .A1(\MR_int[2][16] ), .A2(n956), .ZN(n590) );
  NAND2_X1 U739 ( .A1(\MR_int[2][20] ), .A2(n968), .ZN(n591) );
  AND2_X1 U740 ( .A1(\ML_int[1][1] ), .A2(n987), .ZN(\ML_int[2][1] ) );
  AND2_X1 U741 ( .A1(\ML_int[1][0] ), .A2(n988), .ZN(\ML_int[2][0] ) );
  NAND2_X1 U742 ( .A1(n312), .A2(n313), .ZN(n460) );
  OR2_X1 U743 ( .A1(n684), .A2(n759), .ZN(n312) );
  NOR2_X1 U744 ( .A1(n947), .A2(\SHMAG[5] ), .ZN(n313) );
  NAND2_X1 U745 ( .A1(n182), .A2(n183), .ZN(n759) );
  INV_X1 U746 ( .A(\MR_int[1][31] ), .ZN(n1031) );
  OR2_X1 U747 ( .A1(n948), .A2(\SHMAG[5] ), .ZN(n208) );
  AND2_X1 U748 ( .A1(n982), .A2(\MR_int[1][30] ), .ZN(\MR_int[2][30] ) );
  NAND2_X1 U749 ( .A1(n420), .A2(n419), .ZN(\ML_int[4][28] ) );
  NAND2_X1 U750 ( .A1(n253), .A2(n996), .ZN(n420) );
  NAND2_X1 U751 ( .A1(\ML_int[3][28] ), .A2(n1007), .ZN(n419) );
  NAND2_X1 U752 ( .A1(n418), .A2(n417), .ZN(\ML_int[3][28] ) );
  NAND2_X1 U753 ( .A1(n459), .A2(n458), .ZN(\ML_int[2][21] ) );
  NAND2_X1 U754 ( .A1(\ML_int[1][21] ), .A2(n986), .ZN(n458) );
  NAND2_X1 U755 ( .A1(n413), .A2(n414), .ZN(\ML_int[2][29] ) );
  NAND2_X1 U756 ( .A1(n424), .A2(n971), .ZN(n413) );
  NAND2_X1 U757 ( .A1(\ML_int[1][29] ), .A2(n988), .ZN(n414) );
  NAND2_X1 U758 ( .A1(n494), .A2(net61053), .ZN(\ML_int[4][30] ) );
  NAND2_X1 U759 ( .A1(\ML_int[3][22] ), .A2(n994), .ZN(net61053) );
  NAND2_X1 U760 ( .A1(\ML_int[3][30] ), .A2(n1008), .ZN(n494) );
  NAND2_X1 U761 ( .A1(n135), .A2(n136), .ZN(\MR_int[3][1] ) );
  NAND2_X1 U762 ( .A1(\MR_int[2][1] ), .A2(n957), .ZN(n136) );
  NAND2_X1 U763 ( .A1(\MR_int[2][5] ), .A2(n968), .ZN(n135) );
  NAND2_X1 U764 ( .A1(n144), .A2(n145), .ZN(\ML_int[4][26] ) );
  NAND2_X1 U765 ( .A1(\ML_int[3][18] ), .A2(n995), .ZN(n145) );
  NAND2_X1 U766 ( .A1(\ML_int[3][26] ), .A2(n1008), .ZN(n144) );
  AND2_X1 U767 ( .A1(net61465), .A2(n90), .ZN(n173) );
  NAND2_X1 U769 ( .A1(n380), .A2(n381), .ZN(\MR_int[2][6] ) );
  NAND2_X1 U770 ( .A1(\MR_int[1][6] ), .A2(n978), .ZN(n380) );
  NAND2_X1 U771 ( .A1(\MR_int[1][8] ), .A2(n986), .ZN(n381) );
  NAND2_X1 U772 ( .A1(n696), .A2(n212), .ZN(B[3]) );
  NAND2_X1 U773 ( .A1(n677), .A2(n340), .ZN(B[4]) );
  NAND2_X1 U774 ( .A1(n499), .A2(n500), .ZN(B[8]) );
  NAND2_X1 U775 ( .A1(n443), .A2(n442), .ZN(B[20]) );
  NAND2_X1 U776 ( .A1(n568), .A2(n569), .ZN(B[14]) );
  NAND2_X1 U778 ( .A1(n527), .A2(n526), .ZN(B[24]) );
  NAND2_X1 U779 ( .A1(net61046), .A2(n495), .ZN(B[22]) );
  NAND2_X1 U780 ( .A1(n436), .A2(n435), .ZN(B[18]) );
  OAI21_X1 U781 ( .B1(n674), .B2(n672), .A(n572), .ZN(B[19]) );
  OR2_X1 U782 ( .A1(n703), .A2(n704), .ZN(n515) );
  OR2_X1 U783 ( .A1(n948), .A2(\SHMAG[5] ), .ZN(n704) );
  NAND2_X1 U784 ( .A1(\MR_int[4][24] ), .A2(n1017), .ZN(n703) );
  AND2_X1 U785 ( .A1(\MR_int[3][24] ), .A2(n998), .ZN(\MR_int[4][24] ) );
  NAND2_X1 U786 ( .A1(n311), .A2(n310), .ZN(\ML_int[2][22] ) );
  NAND2_X1 U787 ( .A1(\ML_int[1][20] ), .A2(n978), .ZN(n310) );
  NAND2_X1 U788 ( .A1(\ML_int[1][22] ), .A2(n986), .ZN(n311) );
  BUF_X1 U789 ( .A(\temp_int_SH[1] ), .Z(n984) );
  BUF_X1 U790 ( .A(\temp_int_SH[1] ), .Z(n983) );
  NAND2_X1 U791 ( .A1(\ML_int[2][13] ), .A2(n722), .ZN(n356) );
  AND2_X1 U792 ( .A1(n968), .A2(n1007), .ZN(n722) );
  NAND2_X1 U793 ( .A1(n576), .A2(n577), .ZN(B[2]) );
  NAND2_X1 U794 ( .A1(n529), .A2(n528), .ZN(B[30]) );
  NAND2_X1 U795 ( .A1(n150), .A2(n151), .ZN(\ML_int[3][31] ) );
  NAND2_X1 U796 ( .A1(n250), .A2(n958), .ZN(n150) );
  NAND2_X1 U797 ( .A1(\ML_int[2][31] ), .A2(n968), .ZN(n151) );
  BUF_X1 U798 ( .A(\temp_int_SH[2] ), .Z(n965) );
  BUF_X1 U799 ( .A(\temp_int_SH[2] ), .Z(n966) );
  BUF_X1 U800 ( .A(\temp_int_SH[3] ), .Z(n1005) );
  BUF_X1 U801 ( .A(\temp_int_SH[3] ), .Z(n1006) );
  BUF_X1 U802 ( .A(\temp_int_SH[1] ), .Z(n985) );
  NAND2_X1 U803 ( .A1(SH[5]), .A2(net141507), .ZN(n92) );
  NOR3_X1 U804 ( .A1(n761), .A2(n762), .A3(n763), .ZN(n109) );
  OR2_X1 U805 ( .A1(SH[27]), .A2(SH[26]), .ZN(n761) );
  NAND2_X1 U806 ( .A1(n1047), .A2(n1049), .ZN(n762) );
  NAND2_X1 U807 ( .A1(n1048), .A2(n1050), .ZN(n763) );
  NAND2_X1 U808 ( .A1(net60578), .A2(SH[31]), .ZN(net141507) );
  NAND4_X1 U809 ( .A1(SH[11]), .A2(SH[12]), .A3(SH[13]), .A4(SH[10]), .ZN(
        net60750) );
  NOR2_X1 U810 ( .A1(n1051), .A2(n1032), .ZN(\MR_int[1][31] ) );
  INV_X1 U811 ( .A(A[31]), .ZN(n1051) );
  INV_X1 U812 ( .A(SH[31]), .ZN(n1046) );
  NAND2_X1 U813 ( .A1(n97), .A2(SH[31]), .ZN(n91) );
  NAND4_X1 U814 ( .A1(n101), .A2(n98), .A3(n99), .A4(n100), .ZN(n97) );
  AND2_X1 U815 ( .A1(net60450), .A2(n104), .ZN(n99) );
  NOR2_X1 U816 ( .A1(net60750), .A2(net60751), .ZN(n101) );
  OAI21_X1 U817 ( .B1(n678), .B2(n679), .A(SH[31]), .ZN(n677) );
  AND2_X1 U818 ( .A1(\MR_int[4][5] ), .A2(n205), .ZN(n678) );
  NOR2_X1 U819 ( .A1(n675), .A2(n676), .ZN(n679) );
  NAND2_X1 U820 ( .A1(n127), .A2(n128), .ZN(\MR_int[4][5] ) );
  NAND2_X1 U821 ( .A1(n91), .A2(SH[0]), .ZN(net141444) );
  NAND2_X1 U822 ( .A1(\MR_int[7][20] ), .A2(SH[31]), .ZN(n442) );
  NOR2_X1 U823 ( .A1(n740), .A2(n741), .ZN(\MR_int[7][20] ) );
  AND2_X1 U824 ( .A1(n606), .A2(n607), .ZN(n740) );
  OR2_X1 U825 ( .A1(\SHMAG[5] ), .A2(n1015), .ZN(n741) );
  NAND2_X1 U826 ( .A1(\MR_int[7][24] ), .A2(SH[31]), .ZN(n526) );
  AND2_X1 U827 ( .A1(\MR_int[4][25] ), .A2(n391), .ZN(\MR_int[7][24] ) );
  NAND2_X1 U828 ( .A1(\MR_int[7][30] ), .A2(SH[31]), .ZN(n528) );
  AND2_X1 U829 ( .A1(\MR_int[4][31] ), .A2(n391), .ZN(\MR_int[7][30] ) );
  AND2_X1 U830 ( .A1(n1000), .A2(\MR_int[3][31] ), .ZN(\MR_int[4][31] ) );
  NAND2_X1 U831 ( .A1(\ML_int[1][8] ), .A2(n986), .ZN(n334) );
  NAND2_X1 U832 ( .A1(\MR_int[7][22] ), .A2(SH[31]), .ZN(net61046) );
  NOR3_X1 U833 ( .A1(n1013), .A2(\SHMAG[5] ), .A3(n580), .ZN(\MR_int[7][22] )
         );
  AND2_X1 U834 ( .A1(n602), .A2(n603), .ZN(n580) );
  NAND2_X1 U835 ( .A1(\MR_int[3][23] ), .A2(n997), .ZN(n602) );
  NAND2_X1 U836 ( .A1(SH[4]), .A2(net141507), .ZN(n90) );
  AND3_X1 U837 ( .A1(net60313), .A2(n292), .A3(n291), .ZN(n110) );
  NOR2_X1 U838 ( .A1(SH[6]), .A2(SH[9]), .ZN(n291) );
  NOR2_X1 U839 ( .A1(SH[8]), .A2(SH[7]), .ZN(n292) );
  NOR3_X1 U840 ( .A1(SH[28]), .A2(SH[29]), .A3(SH[30]), .ZN(net60313) );
  NAND2_X1 U841 ( .A1(\ML_int[1][15] ), .A2(n978), .ZN(n302) );
  AND2_X1 U842 ( .A1(n287), .A2(n289), .ZN(n108) );
  NOR3_X1 U843 ( .A1(SH[17]), .A2(SH[18]), .A3(SH[16]), .ZN(n287) );
  NOR3_X1 U844 ( .A1(SH[20]), .A2(SH[21]), .A3(SH[19]), .ZN(n289) );
  NAND2_X1 U845 ( .A1(net61724), .A2(n354), .ZN(\MR_int[2][20] ) );
  NAND2_X1 U846 ( .A1(\MR_int[1][20] ), .A2(n979), .ZN(net61724) );
  NAND2_X1 U847 ( .A1(n186), .A2(n986), .ZN(n354) );
  NAND2_X1 U848 ( .A1(n560), .A2(n561), .ZN(\MR_int[2][22] ) );
  NAND2_X1 U849 ( .A1(\MR_int[1][22] ), .A2(n979), .ZN(n561) );
  NAND2_X1 U850 ( .A1(\MR_int[1][24] ), .A2(n986), .ZN(n560) );
  AND2_X1 U851 ( .A1(n290), .A2(n288), .ZN(n107) );
  NOR3_X1 U852 ( .A1(SH[14]), .A2(SH[15]), .A3(SH[13]), .ZN(n290) );
  NOR3_X1 U853 ( .A1(SH[11]), .A2(SH[12]), .A3(SH[10]), .ZN(n288) );
  NAND2_X1 U854 ( .A1(\ML_int[2][28] ), .A2(n967), .ZN(n417) );
  NAND2_X1 U855 ( .A1(n91), .A2(SH[0]), .ZN(n96) );
  NAND2_X1 U856 ( .A1(\MR_int[1][29] ), .A2(n979), .ZN(n597) );
  NAND2_X1 U857 ( .A1(n732), .A2(n979), .ZN(n571) );
  NAND2_X1 U858 ( .A1(n89), .A2(n95), .ZN(\temp_int_SH[1] ) );
  NAND2_X1 U859 ( .A1(SH[1]), .A2(net60576), .ZN(n95) );
  NAND2_X1 U860 ( .A1(net60578), .A2(SH[31]), .ZN(net60576) );
  NAND2_X1 U861 ( .A1(net61465), .A2(n260), .ZN(\temp_int_SH[2] ) );
  NAND2_X1 U862 ( .A1(SH[2]), .A2(net141507), .ZN(n260) );
  NAND2_X1 U863 ( .A1(net61465), .A2(n717), .ZN(\temp_int_SH[3] ) );
  NAND2_X1 U864 ( .A1(SH[3]), .A2(net141507), .ZN(n717) );
  AND2_X1 U865 ( .A1(n1032), .A2(A[0]), .ZN(\ML_int[1][0] ) );
  AND3_X1 U866 ( .A1(SH[24]), .A2(SH[25]), .A3(SH[23]), .ZN(n104) );
  AND3_X1 U867 ( .A1(SH[28]), .A2(SH[26]), .A3(SH[27]), .ZN(net60450) );
  NAND2_X1 U868 ( .A1(n563), .A2(n562), .ZN(\MR_int[2][26] ) );
  NAND2_X1 U869 ( .A1(\MR_int[1][26] ), .A2(n980), .ZN(n562) );
  NAND2_X1 U870 ( .A1(\MR_int[1][28] ), .A2(n986), .ZN(n563) );
  OR2_X1 U871 ( .A1(n267), .A2(SH[31]), .ZN(n500) );
  NAND2_X1 U872 ( .A1(\ML_int[4][8] ), .A2(n622), .ZN(n267) );
  NAND2_X1 U873 ( .A1(n490), .A2(n491), .ZN(\ML_int[4][8] ) );
  NAND2_X1 U874 ( .A1(\ML_int[3][8] ), .A2(n1009), .ZN(n490) );
  INV_X1 U875 ( .A(SH[22]), .ZN(n1050) );
  INV_X1 U876 ( .A(SH[23]), .ZN(n1049) );
  INV_X1 U877 ( .A(SH[25]), .ZN(n1047) );
  INV_X1 U878 ( .A(SH[24]), .ZN(n1048) );
endmodule


module SHIFTER_M32_N5_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n86, n87, n88, n89, n90, n91, n92, n93, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201,
         n202, n203, n204, n205, n206, n208, n209, n210, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n240, n241, n242, n243, n244, n245, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n260, n263, n265,
         n266, n268, n272, n273, n279, n280, n283, n286, n287, n290, n291,
         n294, n295, n298, n299, n302, n303, n305, n306, n309, n310, n314,
         n315, n316, n317, n318, n321, n322, n325, n326, n327, n329, n330,
         n331, n332, n334, n335, n336, n337, n338, n341, n342, n343, n344,
         n347, n348, n350, n351, n352, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n371, n372,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n385,
         n387, n388, n424, n477, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n570, n571, n572,
         n573, n574, n575, n576, n577, n581, n586, n587, n591, n592, n600,
         n601, n602, n605, n606, n607, n610, n612, n614, n615, n616, n648,
         n668, n699, n700, n701, n702, n703, n763, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974;

  NAND3_X1 U93 ( .A1(n101), .A2(n927), .A3(n102), .ZN(n100) );
  MUX2_X1 U96 ( .A(n109), .B(n110), .S(n111), .Z(n108) );
  MUX2_X1 U98 ( .A(n115), .B(n116), .S(n111), .Z(n114) );
  MUX2_X1 U100 ( .A(n119), .B(n120), .S(n111), .Z(n118) );
  MUX2_X1 U102 ( .A(n123), .B(n124), .S(n111), .Z(n122) );
  MUX2_X1 U104 ( .A(n127), .B(n128), .S(n111), .Z(n126) );
  MUX2_X1 U106 ( .A(n577), .B(n131), .S(n111), .Z(n129) );
  NAND3_X1 U109 ( .A1(n136), .A2(n137), .A3(n132), .ZN(n135) );
  NAND3_X1 U132 ( .A1(n101), .A2(n927), .A3(n170), .ZN(n177) );
  MUX2_X1 U141 ( .A(n182), .B(n183), .S(n111), .Z(n181) );
  NAND3_X1 U197 ( .A1(n136), .A2(n137), .A3(n206), .ZN(n208) );
  MUX2_X1 U244 ( .A(n189), .B(n190), .S(n111), .Z(n227) );
  NAND3_X1 U23 ( .A1(n290), .A2(n291), .A3(n204), .ZN(n263) );
  NAND3_X1 U46 ( .A1(n351), .A2(n350), .A3(n197), .ZN(n142) );
  NAND3_X1 U59 ( .A1(n279), .A2(n280), .A3(n212), .ZN(n162) );
  NAND3_X1 U71 ( .A1(n286), .A2(n287), .A3(n198), .ZN(n144) );
  NAND3_X1 U76 ( .A1(n290), .A2(n291), .A3(n204), .ZN(n149) );
  NAND3_X1 U81 ( .A1(n294), .A2(n295), .A3(n233), .ZN(n152) );
  NAND3_X1 U86 ( .A1(n298), .A2(n299), .A3(n225), .ZN(n176) );
  NAND3_X1 U94 ( .A1(n302), .A2(n303), .A3(n236), .ZN(n158) );
  NAND3_X1 U107 ( .A1(n305), .A2(n306), .A3(n199), .ZN(n148) );
  NAND3_X1 U122 ( .A1(n314), .A2(n315), .A3(n232), .ZN(n157) );
  NAND3_X1 U130 ( .A1(n224), .A2(n338), .A3(n337), .ZN(n321) );
  NAND3_X1 U138 ( .A1(n325), .A2(n326), .A3(n203), .ZN(n145) );
  NAND3_X1 U154 ( .A1(n337), .A2(n338), .A3(n224), .ZN(n172) );
  NAND3_X1 U170 ( .A1(n347), .A2(n348), .A3(n223), .ZN(n169) );
  NAND3_X1 U182 ( .A1(n358), .A2(n359), .A3(n217), .ZN(n164) );
  NAND3_X1 U190 ( .A1(n365), .A2(n366), .A3(n216), .ZN(n167) );
  NAND3_X1 U193 ( .A1(n367), .A2(n368), .A3(n235), .ZN(n150) );
  NAND3_X1 U200 ( .A1(n371), .A2(n372), .A3(n202), .ZN(n141) );
  NAND3_X1 U208 ( .A1(n215), .A2(n380), .A3(n379), .ZN(n163) );
  NAND3_X1 U373 ( .A1(SH[15]), .A2(SH[14]), .A3(SH[16]), .ZN(n506) );
  NAND3_X1 U22 ( .A1(n317), .A2(n318), .A3(n221), .ZN(n571) );
  MUX2_X1 U34 ( .A(n160), .B(n159), .S(n196), .Z(n136) );
  NAND3_X1 U44 ( .A1(n336), .A2(n335), .A3(n230), .ZN(n154) );
  NAND3_X1 U45 ( .A1(n209), .A2(n343), .A3(n342), .ZN(n159) );
  NAND3_X1 U47 ( .A1(n364), .A2(n363), .A3(n362), .ZN(n648) );
  NAND3_X1 U52 ( .A1(n331), .A2(n332), .A3(n210), .ZN(n586) );
  NAND3_X1 U53 ( .A1(n294), .A2(n295), .A3(n233), .ZN(n587) );
  NAND3_X1 U60 ( .A1(n358), .A2(n359), .A3(n217), .ZN(n592) );
  NAND3_X1 U70 ( .A1(n279), .A2(n280), .A3(n212), .ZN(n600) );
  NAND3_X1 U73 ( .A1(n215), .A2(n380), .A3(n379), .ZN(n602) );
  NAND3_X1 U309 ( .A1(n354), .A2(n355), .A3(n226), .ZN(n173) );
  NAND3_X1 U311 ( .A1(n317), .A2(n318), .A3(n221), .ZN(n168) );
  NAND3_X1 U317 ( .A1(n331), .A2(n332), .A3(n210), .ZN(n166) );
  MUX2_X1 U128 ( .A(n142), .B(n143), .S(n196), .Z(n101) );
  AOI222_X1 U3 ( .A1(n912), .A2(A[1]), .B1(n915), .B2(A[0]), .C1(n935), .C2(
        A[2]), .ZN(n106) );
  BUF_X1 U4 ( .A(n926), .Z(n899) );
  BUF_X1 U5 ( .A(n926), .Z(n898) );
  BUF_X1 U6 ( .A(n926), .Z(n900) );
  INV_X1 U7 ( .A(n132), .ZN(n916) );
  BUF_X1 U8 ( .A(n928), .Z(n902) );
  BUF_X1 U9 ( .A(n931), .Z(n904) );
  BUF_X1 U10 ( .A(n928), .Z(n901) );
  BUF_X1 U11 ( .A(n931), .Z(n905) );
  INV_X1 U12 ( .A(n170), .ZN(n918) );
  BUF_X1 U13 ( .A(n931), .Z(n906) );
  NAND2_X1 U14 ( .A1(n132), .A2(n898), .ZN(n112) );
  NAND2_X1 U15 ( .A1(n170), .A2(n901), .ZN(n179) );
  INV_X1 U16 ( .A(n614), .ZN(n926) );
  BUF_X1 U17 ( .A(n928), .Z(n903) );
  AOI222_X1 U18 ( .A1(n600), .A2(n905), .B1(n934), .B2(n908), .C1(n586), .C2(
        n901), .ZN(n133) );
  INV_X1 U19 ( .A(n102), .ZN(n919) );
  NOR2_X1 U20 ( .A1(n107), .A2(n921), .ZN(n132) );
  AOI22_X1 U21 ( .A1(n587), .A2(n901), .B1(n572), .B2(n905), .ZN(n91) );
  AOI22_X1 U24 ( .A1(n571), .A2(n898), .B1(n938), .B2(n908), .ZN(n140) );
  INV_X1 U25 ( .A(n206), .ZN(n917) );
  BUF_X1 U26 ( .A(n272), .Z(n914) );
  BUF_X1 U27 ( .A(n272), .Z(n913) );
  BUF_X1 U28 ( .A(n387), .Z(n907) );
  BUF_X1 U29 ( .A(n385), .Z(n911) );
  BUF_X1 U30 ( .A(n385), .Z(n910) );
  BUF_X1 U31 ( .A(n387), .Z(n908) );
  BUF_X1 U32 ( .A(n272), .Z(n915) );
  NOR2_X1 U33 ( .A1(n113), .A2(n921), .ZN(n170) );
  BUF_X1 U35 ( .A(n385), .Z(n912) );
  NOR3_X1 U36 ( .A1(n376), .A2(n375), .A3(n374), .ZN(n341) );
  NOR3_X1 U37 ( .A1(n381), .A2(n382), .A3(n923), .ZN(n316) );
  NOR3_X1 U38 ( .A1(n329), .A2(n330), .A3(n925), .ZN(n92) );
  INV_X1 U39 ( .A(n165), .ZN(n925) );
  AOI22_X1 U40 ( .A1(n899), .A2(n934), .B1(n902), .B2(n602), .ZN(n192) );
  BUF_X1 U41 ( .A(n387), .Z(n909) );
  NAND2_X1 U42 ( .A1(n102), .A2(n901), .ZN(n104) );
  NAND2_X1 U43 ( .A1(n206), .A2(n898), .ZN(n191) );
  INV_X1 U48 ( .A(n273), .ZN(n939) );
  INV_X1 U49 ( .A(n572), .ZN(n936) );
  INV_X1 U50 ( .A(n334), .ZN(n935) );
  OR2_X1 U51 ( .A1(n932), .A2(n927), .ZN(n614) );
  INV_X1 U54 ( .A(n615), .ZN(n928) );
  INV_X1 U55 ( .A(n763), .ZN(n931) );
  AND2_X1 U56 ( .A1(n136), .A2(n927), .ZN(n376) );
  AND3_X1 U57 ( .A1(n499), .A2(n500), .A3(n184), .ZN(n110) );
  NAND2_X1 U58 ( .A1(n586), .A2(n907), .ZN(n499) );
  NAND2_X1 U61 ( .A1(n602), .A2(n904), .ZN(n500) );
  AOI22_X1 U62 ( .A1(n600), .A2(n898), .B1(n902), .B2(n592), .ZN(n184) );
  INV_X1 U63 ( .A(n143), .ZN(n937) );
  INV_X1 U64 ( .A(n160), .ZN(n940) );
  AND3_X1 U65 ( .A1(n192), .A2(n930), .A3(n922), .ZN(n352) );
  INV_X1 U66 ( .A(n378), .ZN(n930) );
  INV_X1 U67 ( .A(n377), .ZN(n922) );
  OAI221_X1 U68 ( .B1(n98), .B2(n917), .C1(n99), .C2(n916), .A(n100), .ZN(B[5]) );
  OAI222_X1 U69 ( .A1(n95), .A2(n916), .B1(n96), .B2(n917), .C1(n97), .C2(n919), .ZN(B[6]) );
  OAI221_X1 U72 ( .B1(n919), .B2(n929), .C1(n917), .C2(n93), .A(n570), .ZN(
        B[7]) );
  OAI222_X1 U74 ( .A1(n86), .A2(n916), .B1(n87), .B2(n917), .C1(n88), .C2(n919), .ZN(B[9]) );
  OAI22_X1 U75 ( .A1(n940), .A2(n112), .B1(n113), .B2(n114), .ZN(B[31]) );
  OAI222_X1 U77 ( .A1(n138), .A2(n916), .B1(n140), .B2(n917), .C1(n139), .C2(
        n919), .ZN(B[10]) );
  OAI222_X1 U78 ( .A1(n92), .A2(n919), .B1(n929), .B2(n918), .C1(n93), .C2(
        n916), .ZN(B[23]) );
  OAI222_X1 U79 ( .A1(n127), .A2(n916), .B1(n125), .B2(n191), .C1(n322), .C2(
        n919), .ZN(B[13]) );
  OAI222_X1 U80 ( .A1(n577), .A2(n916), .B1(n942), .B2(n191), .C1(n131), .C2(
        n919), .ZN(B[12]) );
  OAI222_X1 U82 ( .A1(n388), .A2(n916), .B1(n940), .B2(n191), .C1(n352), .C2(
        n919), .ZN(B[15]) );
  OAI222_X1 U83 ( .A1(n183), .A2(n919), .B1(n937), .B2(n179), .C1(n182), .C2(
        n916), .ZN(B[17]) );
  OAI222_X1 U84 ( .A1(n86), .A2(n919), .B1(n88), .B2(n918), .C1(n87), .C2(n916), .ZN(B[25]) );
  OAI222_X1 U85 ( .A1(n138), .A2(n919), .B1(n139), .B2(n918), .C1(n140), .C2(
        n916), .ZN(B[26]) );
  OR2_X1 U87 ( .A1(n268), .A2(n916), .ZN(n570) );
  AND2_X1 U88 ( .A1(n165), .A2(n612), .ZN(n268) );
  NOR2_X1 U89 ( .A1(n330), .A2(n329), .ZN(n612) );
  OAI221_X1 U90 ( .B1(n133), .B2(n918), .C1(n134), .C2(n919), .A(n135), .ZN(
        B[27]) );
  OAI221_X1 U91 ( .B1(n134), .B2(n916), .C1(n133), .C2(n919), .A(n208), .ZN(
        B[11]) );
  OAI221_X1 U92 ( .B1(n99), .B2(n919), .C1(n98), .C2(n916), .A(n177), .ZN(
        B[21]) );
  OAI22_X1 U95 ( .A1(n937), .A2(n104), .B1(n107), .B2(n181), .ZN(B[1]) );
  OAI22_X1 U97 ( .A1(n942), .A2(n112), .B1(n113), .B2(n129), .ZN(B[28]) );
  AOI222_X1 U99 ( .A1(n938), .A2(n906), .B1(n571), .B2(n908), .C1(n169), .C2(
        n898), .ZN(n96) );
  AOI222_X1 U101 ( .A1(n142), .A2(n906), .B1(n909), .B2(n143), .C1(n144), .C2(
        n901), .ZN(n88) );
  AOI222_X1 U103 ( .A1(n171), .A2(n905), .B1(n933), .B2(n908), .C1(n175), .C2(
        n901), .ZN(n139) );
  AOI222_X1 U105 ( .A1(n159), .A2(n908), .B1(n906), .B2(n160), .C1(n161), .C2(
        n898), .ZN(n93) );
  AOI222_X1 U108 ( .A1(n151), .A2(n905), .B1(n150), .B2(n908), .C1(n158), .C2(
        n898), .ZN(n103) );
  AOI222_X1 U110 ( .A1(n648), .A2(n905), .B1(n141), .B2(n908), .C1(n263), .C2(
        n898), .ZN(n98) );
  AOI222_X1 U111 ( .A1(n148), .A2(n901), .B1(n144), .B2(n905), .C1(n137), .C2(
        n101), .ZN(n322) );
  AOI221_X1 U112 ( .B1(n152), .B2(n909), .C1(n157), .C2(n904), .A(n668), .ZN(
        n190) );
  OAI22_X1 U113 ( .A1(n266), .A2(n615), .B1(n936), .B2(n614), .ZN(n668) );
  NAND2_X1 U114 ( .A1(n240), .A2(n943), .ZN(n616) );
  OAI221_X1 U115 ( .B1(n273), .B2(n974), .C1(n334), .C2(n972), .A(n231), .ZN(
        n572) );
  AOI221_X1 U116 ( .B1(n167), .B2(n909), .C1(n161), .C2(n904), .A(n924), .ZN(
        n388) );
  NAND2_X1 U117 ( .A1(n943), .A2(n240), .ZN(n273) );
  OR2_X1 U118 ( .A1(n240), .A2(n943), .ZN(n334) );
  OR2_X1 U119 ( .A1(n240), .A2(n943), .ZN(n591) );
  OAI221_X1 U120 ( .B1(n273), .B2(n974), .C1(n334), .C2(n972), .A(n231), .ZN(
        n153) );
  NOR2_X1 U121 ( .A1(n113), .A2(n111), .ZN(n102) );
  AOI22_X1 U123 ( .A1(n171), .A2(n901), .B1(n933), .B2(n905), .ZN(n97) );
  AOI22_X1 U124 ( .A1(n150), .A2(n898), .B1(n151), .B2(n908), .ZN(n90) );
  AOI22_X1 U125 ( .A1(n141), .A2(n898), .B1(n648), .B2(n908), .ZN(n87) );
  NAND2_X1 U126 ( .A1(n218), .A2(n920), .ZN(n107) );
  AOI22_X1 U127 ( .A1(n899), .A2(n586), .B1(n902), .B2(n167), .ZN(n165) );
  NOR2_X1 U129 ( .A1(n107), .A2(n111), .ZN(n206) );
  NOR2_X1 U131 ( .A1(n273), .A2(n944), .ZN(n160) );
  OR2_X1 U133 ( .A1(n920), .A2(n218), .ZN(n113) );
  NOR2_X1 U134 ( .A1(n974), .A2(n334), .ZN(n143) );
  NOR2_X1 U135 ( .A1(n107), .A2(n227), .ZN(B[0]) );
  INV_X1 U136 ( .A(n383), .ZN(n943) );
  INV_X1 U137 ( .A(n137), .ZN(n927) );
  INV_X1 U139 ( .A(n106), .ZN(n934) );
  NOR2_X1 U140 ( .A1(n240), .A2(n383), .ZN(n272) );
  OR2_X1 U142 ( .A1(n196), .A2(n137), .ZN(n615) );
  NOR2_X1 U143 ( .A1(n196), .A2(n927), .ZN(n387) );
  NOR2_X1 U144 ( .A1(n424), .A2(n576), .ZN(n577) );
  NAND2_X1 U145 ( .A1(n574), .A2(n575), .ZN(n576) );
  OAI22_X1 U146 ( .A1(n615), .A2(n265), .B1(n614), .B2(n266), .ZN(n424) );
  NAND2_X1 U147 ( .A1(n158), .A2(n904), .ZN(n575) );
  INV_X1 U148 ( .A(n117), .ZN(n938) );
  NAND2_X1 U149 ( .A1(n155), .A2(n908), .ZN(n574) );
  INV_X1 U150 ( .A(n151), .ZN(n942) );
  INV_X1 U151 ( .A(n121), .ZN(n933) );
  INV_X1 U152 ( .A(n111), .ZN(n921) );
  AND2_X1 U153 ( .A1(n240), .A2(n383), .ZN(n385) );
  AND3_X1 U155 ( .A1(n481), .A2(n482), .A3(n180), .ZN(n105) );
  NAND2_X1 U156 ( .A1(n154), .A2(n905), .ZN(n482) );
  NAND2_X1 U157 ( .A1(n157), .A2(n908), .ZN(n481) );
  AOI22_X1 U158 ( .A1(n899), .A2(n587), .B1(n155), .B2(n901), .ZN(n180) );
  AND3_X1 U159 ( .A1(n336), .A2(n335), .A3(n230), .ZN(n266) );
  AND3_X1 U160 ( .A1(n483), .A2(n484), .A3(n178), .ZN(n99) );
  NAND2_X1 U161 ( .A1(n145), .A2(n905), .ZN(n484) );
  NAND2_X1 U162 ( .A1(n148), .A2(n907), .ZN(n483) );
  AOI22_X1 U163 ( .A1(n899), .A2(n144), .B1(n902), .B2(n146), .ZN(n178) );
  AND3_X1 U164 ( .A1(n699), .A2(n700), .A3(n213), .ZN(n134) );
  NAND2_X1 U165 ( .A1(n592), .A2(n907), .ZN(n699) );
  NAND2_X1 U166 ( .A1(n167), .A2(n904), .ZN(n700) );
  AOI22_X1 U167 ( .A1(n899), .A2(n602), .B1(n601), .B2(n901), .ZN(n213) );
  AND3_X1 U168 ( .A1(n485), .A2(n486), .A3(n147), .ZN(n86) );
  NAND2_X1 U169 ( .A1(n145), .A2(n907), .ZN(n485) );
  NAND2_X1 U171 ( .A1(n146), .A2(n905), .ZN(n486) );
  AOI22_X1 U172 ( .A1(n899), .A2(n148), .B1(n902), .B2(n149), .ZN(n147) );
  AND3_X1 U173 ( .A1(n489), .A2(n490), .A3(n156), .ZN(n89) );
  NAND2_X1 U174 ( .A1(n154), .A2(n907), .ZN(n489) );
  NAND2_X1 U175 ( .A1(n155), .A2(n905), .ZN(n490) );
  AOI22_X1 U176 ( .A1(n899), .A2(n157), .B1(n902), .B2(n158), .ZN(n156) );
  AND3_X1 U177 ( .A1(n487), .A2(n488), .A3(n174), .ZN(n95) );
  NAND2_X1 U178 ( .A1(n321), .A2(n907), .ZN(n487) );
  NAND2_X1 U179 ( .A1(n173), .A2(n905), .ZN(n488) );
  AOI22_X1 U180 ( .A1(n175), .A2(n898), .B1(n902), .B2(n176), .ZN(n174) );
  AND3_X1 U181 ( .A1(n491), .A2(n492), .A3(n222), .ZN(n138) );
  NAND2_X1 U183 ( .A1(n176), .A2(n904), .ZN(n492) );
  NAND2_X1 U184 ( .A1(n173), .A2(n907), .ZN(n491) );
  AOI22_X1 U185 ( .A1(n899), .A2(n321), .B1(n902), .B2(n169), .ZN(n222) );
  AND3_X1 U186 ( .A1(n362), .A2(n363), .A3(n364), .ZN(n125) );
  NOR3_X1 U187 ( .A1(n381), .A2(n382), .A3(n923), .ZN(n119) );
  AND2_X1 U188 ( .A1(n192), .A2(n310), .ZN(n116) );
  NOR3_X1 U189 ( .A1(n356), .A2(n357), .A3(n924), .ZN(n115) );
  NOR2_X1 U191 ( .A1(n378), .A2(n377), .ZN(n310) );
  AND2_X1 U192 ( .A1(n167), .A2(n900), .ZN(n374) );
  AND2_X1 U194 ( .A1(n601), .A2(n909), .ZN(n375) );
  AND2_X1 U195 ( .A1(n169), .A2(n906), .ZN(n382) );
  AND2_X1 U196 ( .A1(n176), .A2(n909), .ZN(n381) );
  NOR3_X1 U198 ( .A1(n605), .A2(n606), .A3(n607), .ZN(n128) );
  AND2_X1 U199 ( .A1(n137), .A2(n101), .ZN(n607) );
  AND2_X1 U201 ( .A1(n148), .A2(n903), .ZN(n605) );
  NOR3_X1 U202 ( .A1(n376), .A2(n375), .A3(n374), .ZN(n109) );
  AND2_X1 U203 ( .A1(n164), .A2(n906), .ZN(n330) );
  AND2_X1 U204 ( .A1(n163), .A2(n909), .ZN(n329) );
  AND2_X1 U205 ( .A1(n162), .A2(n909), .ZN(n377) );
  AND2_X1 U206 ( .A1(n166), .A2(n906), .ZN(n378) );
  INV_X1 U207 ( .A(n193), .ZN(n924) );
  AOI22_X1 U209 ( .A1(n899), .A2(n592), .B1(n902), .B2(n159), .ZN(n193) );
  INV_X1 U210 ( .A(n195), .ZN(n923) );
  AOI22_X1 U211 ( .A1(n899), .A2(n173), .B1(n902), .B2(n168), .ZN(n195) );
  AND3_X1 U212 ( .A1(n493), .A2(n494), .A3(n185), .ZN(n123) );
  NAND2_X1 U213 ( .A1(n168), .A2(n904), .ZN(n494) );
  NAND2_X1 U214 ( .A1(n169), .A2(n907), .ZN(n493) );
  AOI22_X1 U215 ( .A1(n900), .A2(n176), .B1(n902), .B2(n938), .ZN(n185) );
  INV_X1 U216 ( .A(n581), .ZN(n929) );
  OAI22_X1 U217 ( .A1(n615), .A2(n941), .B1(n106), .B2(n763), .ZN(n581) );
  INV_X1 U218 ( .A(n600), .ZN(n941) );
  AND3_X1 U219 ( .A1(n701), .A2(n702), .A3(n703), .ZN(n131) );
  NAND2_X1 U220 ( .A1(n152), .A2(n904), .ZN(n701) );
  NAND2_X1 U221 ( .A1(n153), .A2(n907), .ZN(n702) );
  NAND2_X1 U222 ( .A1(n157), .A2(n901), .ZN(n703) );
  AND3_X1 U223 ( .A1(n186), .A2(n260), .A3(n477), .ZN(n124) );
  NAND2_X1 U224 ( .A1(n172), .A2(n904), .ZN(n260) );
  NAND2_X1 U225 ( .A1(n175), .A2(n907), .ZN(n477) );
  AOI22_X1 U226 ( .A1(n900), .A2(n171), .B1(n902), .B2(n173), .ZN(n186) );
  AND3_X1 U227 ( .A1(n495), .A2(n496), .A3(n201), .ZN(n127) );
  NAND2_X1 U228 ( .A1(n149), .A2(n904), .ZN(n496) );
  NAND2_X1 U229 ( .A1(n146), .A2(n907), .ZN(n495) );
  AOI22_X1 U230 ( .A1(n900), .A2(n145), .B1(n903), .B2(n141), .ZN(n201) );
  AND3_X1 U231 ( .A1(n497), .A2(n498), .A3(n188), .ZN(n183) );
  NAND2_X1 U232 ( .A1(n144), .A2(n907), .ZN(n497) );
  NAND2_X1 U233 ( .A1(n148), .A2(n904), .ZN(n498) );
  AOI22_X1 U234 ( .A1(n899), .A2(n142), .B1(n903), .B2(n145), .ZN(n188) );
  AND3_X1 U235 ( .A1(n501), .A2(n502), .A3(n234), .ZN(n189) );
  NAND2_X1 U236 ( .A1(n155), .A2(n898), .ZN(n501) );
  NAND2_X1 U237 ( .A1(n151), .A2(n901), .ZN(n502) );
  AOI22_X1 U238 ( .A1(n909), .A2(n158), .B1(n906), .B2(n150), .ZN(n234) );
  OR2_X1 U239 ( .A1(n932), .A2(n137), .ZN(n763) );
  AND3_X1 U240 ( .A1(n503), .A2(n504), .A3(n194), .ZN(n120) );
  NAND2_X1 U241 ( .A1(n175), .A2(n904), .ZN(n504) );
  NAND2_X1 U242 ( .A1(n171), .A2(n908), .ZN(n503) );
  AOI22_X1 U243 ( .A1(n899), .A2(n933), .B1(n902), .B2(n172), .ZN(n194) );
  AND3_X1 U245 ( .A1(n367), .A2(n368), .A3(n235), .ZN(n265) );
  INV_X1 U246 ( .A(n196), .ZN(n932) );
  AND2_X1 U247 ( .A1(n327), .A2(n187), .ZN(n182) );
  NOR2_X1 U248 ( .A1(n360), .A2(n361), .ZN(n327) );
  AOI22_X1 U249 ( .A1(n899), .A2(n146), .B1(n902), .B2(n648), .ZN(n187) );
  AND2_X1 U250 ( .A1(n263), .A2(n909), .ZN(n360) );
  AND2_X1 U251 ( .A1(n161), .A2(n906), .ZN(n357) );
  AND2_X1 U252 ( .A1(n144), .A2(n906), .ZN(n606) );
  AND2_X1 U253 ( .A1(n167), .A2(n909), .ZN(n356) );
  AND2_X1 U254 ( .A1(n141), .A2(n906), .ZN(n361) );
  OR2_X1 U255 ( .A1(n616), .A2(n963), .ZN(n335) );
  OR2_X1 U256 ( .A1(n616), .A2(n954), .ZN(n290) );
  OR2_X1 U257 ( .A1(n273), .A2(n964), .ZN(n379) );
  OR2_X1 U258 ( .A1(n273), .A2(n965), .ZN(n337) );
  OR2_X1 U259 ( .A1(n273), .A2(n951), .ZN(n367) );
  OR2_X1 U260 ( .A1(n273), .A2(n972), .ZN(n279) );
  OR2_X1 U261 ( .A1(n273), .A2(n968), .ZN(n331) );
  OR2_X1 U262 ( .A1(n273), .A2(n949), .ZN(n317) );
  OR2_X1 U263 ( .A1(n273), .A2(n971), .ZN(n294) );
  OAI22_X1 U264 ( .A1(n108), .A2(n107), .B1(n104), .B2(n106), .ZN(B[3]) );
  OAI222_X1 U265 ( .A1(n103), .A2(n917), .B1(n936), .B2(n104), .C1(n105), .C2(
        n916), .ZN(B[4]) );
  OAI222_X1 U266 ( .A1(n89), .A2(n916), .B1(n90), .B2(n917), .C1(n91), .C2(
        n919), .ZN(B[8]) );
  OR2_X1 U267 ( .A1(n334), .A2(n961), .ZN(n380) );
  OR2_X1 U268 ( .A1(n334), .A2(n965), .ZN(n332) );
  OR2_X1 U269 ( .A1(n334), .A2(n968), .ZN(n295) );
  OR2_X1 U270 ( .A1(n591), .A2(n957), .ZN(n359) );
  OR2_X1 U271 ( .A1(n591), .A2(n969), .ZN(n280) );
  OR2_X1 U272 ( .A1(n591), .A2(n951), .ZN(n291) );
  OR2_X1 U273 ( .A1(n591), .A2(n962), .ZN(n338) );
  OR2_X1 U274 ( .A1(n948), .A2(n334), .ZN(n368) );
  OAI222_X1 U275 ( .A1(n105), .A2(n919), .B1(n936), .B2(n179), .C1(n103), .C2(
        n916), .ZN(B[20]) );
  OAI222_X1 U276 ( .A1(n316), .A2(n916), .B1(n117), .B2(n191), .C1(n919), .C2(
        n120), .ZN(B[14]) );
  OAI222_X1 U277 ( .A1(n89), .A2(n919), .B1(n91), .B2(n918), .C1(n90), .C2(
        n916), .ZN(B[24]) );
  OAI222_X1 U278 ( .A1(n95), .A2(n919), .B1(n97), .B2(n918), .C1(n96), .C2(
        n916), .ZN(B[22]) );
  OAI222_X1 U279 ( .A1(n124), .A2(n919), .B1(n121), .B2(n179), .C1(n123), .C2(
        n916), .ZN(B[18]) );
  OAI222_X1 U280 ( .A1(n110), .A2(n919), .B1(n106), .B2(n179), .C1(n341), .C2(
        n916), .ZN(B[19]) );
  OAI22_X1 U281 ( .A1(n121), .A2(n104), .B1(n107), .B2(n122), .ZN(B[2]) );
  OAI22_X1 U282 ( .A1(n117), .A2(n112), .B1(n113), .B2(n118), .ZN(B[30]) );
  OAI221_X1 U283 ( .B1(n273), .B2(n958), .C1(n334), .C2(n955), .A(n205), .ZN(
        n146) );
  AOI22_X1 U284 ( .A1(A[18]), .A2(n915), .B1(A[19]), .B2(n912), .ZN(n205) );
  OAI221_X1 U285 ( .B1(n616), .B2(n973), .C1(n591), .C2(n970), .A(n220), .ZN(
        n171) );
  INV_X1 U286 ( .A(A[2]), .ZN(n973) );
  AOI22_X1 U287 ( .A1(A[3]), .A2(n915), .B1(A[4]), .B2(n912), .ZN(n220) );
  OAI221_X1 U288 ( .B1(n273), .B2(n947), .C1(n944), .C2(n591), .A(n237), .ZN(
        n151) );
  AOI22_X1 U289 ( .A1(A[29]), .A2(n915), .B1(n912), .B2(A[30]), .ZN(n237) );
  OAI221_X1 U290 ( .B1(n616), .B2(n969), .C1(n334), .C2(n966), .A(n219), .ZN(
        n175) );
  AOI22_X1 U291 ( .A1(A[7]), .A2(n915), .B1(A[8]), .B2(n912), .ZN(n219) );
  OAI221_X1 U292 ( .B1(n616), .B2(n959), .C1(n334), .C2(n956), .A(n238), .ZN(
        n155) );
  AOI22_X1 U293 ( .A1(A[17]), .A2(n915), .B1(A[18]), .B2(n911), .ZN(n238) );
  OAI221_X1 U294 ( .B1(n616), .B2(n952), .C1(n949), .C2(n334), .A(n573), .ZN(
        n161) );
  AOI22_X1 U295 ( .A1(A[24]), .A2(n914), .B1(A[25]), .B2(n911), .ZN(n573) );
  OR2_X1 U296 ( .A1(n591), .A2(n963), .ZN(n306) );
  OR2_X1 U297 ( .A1(n273), .A2(n966), .ZN(n305) );
  AOI22_X1 U298 ( .A1(A[10]), .A2(n913), .B1(A[11]), .B2(n910), .ZN(n199) );
  OR2_X1 U299 ( .A1(n334), .A2(n967), .ZN(n287) );
  OR2_X1 U300 ( .A1(n616), .A2(n970), .ZN(n286) );
  AOI22_X1 U301 ( .A1(A[6]), .A2(n913), .B1(A[7]), .B2(n910), .ZN(n198) );
  NOR4_X1 U302 ( .A1(n255), .A2(SH[28]), .A3(SH[30]), .A4(SH[29]), .ZN(n254)
         );
  OR4_X1 U303 ( .A1(SH[6]), .A2(SH[7]), .A3(SH[8]), .A4(SH[9]), .ZN(n255) );
  OR2_X1 U304 ( .A1(n591), .A2(n953), .ZN(n366) );
  OR2_X1 U305 ( .A1(n273), .A2(n956), .ZN(n365) );
  AOI22_X1 U306 ( .A1(A[20]), .A2(n913), .B1(A[21]), .B2(n910), .ZN(n216) );
  NOR4_X1 U307 ( .A1(n256), .A2(SH[22]), .A3(SH[24]), .A4(SH[23]), .ZN(n253)
         );
  OR3_X1 U308 ( .A1(SH[26]), .A2(SH[27]), .A3(SH[25]), .ZN(n256) );
  OR2_X1 U310 ( .A1(n334), .A2(n959), .ZN(n326) );
  OR2_X1 U312 ( .A1(n616), .A2(n962), .ZN(n325) );
  AOI22_X1 U313 ( .A1(A[14]), .A2(n913), .B1(A[15]), .B2(n910), .ZN(n203) );
  OR2_X1 U314 ( .A1(n591), .A2(n958), .ZN(n355) );
  OR2_X1 U315 ( .A1(n616), .A2(n961), .ZN(n354) );
  AOI22_X1 U316 ( .A1(A[15]), .A2(n913), .B1(A[16]), .B2(n910), .ZN(n226) );
  OR2_X1 U318 ( .A1(n591), .A2(n952), .ZN(n303) );
  OR2_X1 U319 ( .A1(n616), .A2(n955), .ZN(n302) );
  AOI22_X1 U320 ( .A1(A[21]), .A2(n913), .B1(A[22]), .B2(n910), .ZN(n236) );
  OR2_X1 U321 ( .A1(n591), .A2(n964), .ZN(n315) );
  OR2_X1 U322 ( .A1(n616), .A2(n967), .ZN(n314) );
  AOI22_X1 U323 ( .A1(A[9]), .A2(n913), .B1(A[10]), .B2(n910), .ZN(n232) );
  AOI22_X1 U324 ( .A1(A[30]), .A2(n939), .B1(n915), .B2(A[31]), .ZN(n117) );
  AOI22_X1 U325 ( .A1(n935), .A2(A[1]), .B1(n912), .B2(A[0]), .ZN(n121) );
  OAI221_X1 U326 ( .B1(n616), .B2(n952), .C1(n949), .C2(n334), .A(n214), .ZN(
        n601) );
  AOI22_X1 U327 ( .A1(A[24]), .A2(n913), .B1(A[25]), .B2(n910), .ZN(n214) );
  NAND2_X1 U328 ( .A1(SH[4]), .A2(n228), .ZN(n111) );
  OR2_X1 U329 ( .A1(n334), .A2(n954), .ZN(n299) );
  OR2_X1 U330 ( .A1(n273), .A2(n957), .ZN(n298) );
  AOI22_X1 U331 ( .A1(A[19]), .A2(n913), .B1(A[20]), .B2(n910), .ZN(n225) );
  OR2_X1 U332 ( .A1(n591), .A2(n947), .ZN(n372) );
  OR2_X1 U333 ( .A1(n273), .A2(n950), .ZN(n371) );
  AOI22_X1 U334 ( .A1(A[26]), .A2(n913), .B1(A[27]), .B2(n910), .ZN(n202) );
  OR2_X1 U335 ( .A1(n950), .A2(n334), .ZN(n348) );
  OR2_X1 U336 ( .A1(n273), .A2(n953), .ZN(n347) );
  AOI22_X1 U337 ( .A1(A[23]), .A2(n913), .B1(A[24]), .B2(n910), .ZN(n223) );
  AOI22_X1 U338 ( .A1(A[1]), .A2(n914), .B1(A[2]), .B2(n911), .ZN(n231) );
  NAND2_X1 U339 ( .A1(n344), .A2(SH[0]), .ZN(n240) );
  NAND2_X1 U340 ( .A1(SH[31]), .A2(n283), .ZN(n228) );
  NAND4_X1 U341 ( .A1(n244), .A2(n243), .A3(n245), .A4(n610), .ZN(n283) );
  AND4_X1 U342 ( .A1(n249), .A2(SH[9]), .A3(SH[7]), .A4(SH[8]), .ZN(n610) );
  OR2_X1 U343 ( .A1(n945), .A2(n334), .ZN(n343) );
  OR2_X1 U344 ( .A1(n273), .A2(n948), .ZN(n342) );
  AOI22_X1 U345 ( .A1(A[28]), .A2(n914), .B1(A[29]), .B2(n911), .ZN(n209) );
  OR2_X1 U346 ( .A1(n334), .A2(n971), .ZN(n351) );
  NAND2_X1 U347 ( .A1(n939), .A2(A[1]), .ZN(n350) );
  AOI22_X1 U348 ( .A1(A[2]), .A2(n913), .B1(A[3]), .B2(n910), .ZN(n197) );
  AOI22_X1 U349 ( .A1(n915), .A2(A[25]), .B1(A[26]), .B2(n912), .ZN(n235) );
  NAND2_X1 U350 ( .A1(SH[3]), .A2(n228), .ZN(n137) );
  NAND2_X1 U351 ( .A1(SH[2]), .A2(n228), .ZN(n196) );
  AOI21_X1 U352 ( .B1(n250), .B2(n920), .A(SH[5]), .ZN(n218) );
  NAND4_X1 U353 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(n250) );
  NOR4_X1 U354 ( .A1(n258), .A2(SH[10]), .A3(SH[12]), .A4(SH[11]), .ZN(n251)
         );
  NOR4_X1 U355 ( .A1(n257), .A2(SH[16]), .A3(SH[18]), .A4(SH[17]), .ZN(n252)
         );
  AOI22_X1 U356 ( .A1(A[16]), .A2(n914), .B1(n912), .B2(A[17]), .ZN(n217) );
  AOI22_X1 U357 ( .A1(A[13]), .A2(n914), .B1(A[14]), .B2(n911), .ZN(n230) );
  AOI22_X1 U358 ( .A1(A[4]), .A2(n914), .B1(A[5]), .B2(n911), .ZN(n212) );
  AOI22_X1 U359 ( .A1(A[8]), .A2(n914), .B1(A[9]), .B2(n911), .ZN(n210) );
  AOI22_X1 U360 ( .A1(A[22]), .A2(n914), .B1(A[23]), .B2(n911), .ZN(n204) );
  AOI22_X1 U361 ( .A1(A[27]), .A2(n914), .B1(A[28]), .B2(n911), .ZN(n221) );
  AOI22_X1 U362 ( .A1(A[5]), .A2(n914), .B1(A[6]), .B2(n911), .ZN(n233) );
  AOI22_X1 U363 ( .A1(A[11]), .A2(n914), .B1(A[12]), .B2(n911), .ZN(n224) );
  AOI22_X1 U364 ( .A1(A[12]), .A2(n914), .B1(A[13]), .B2(n911), .ZN(n215) );
  NOR2_X1 U365 ( .A1(n505), .A2(n506), .ZN(n245) );
  NAND4_X1 U366 ( .A1(SH[10]), .A2(SH[12]), .A3(SH[11]), .A4(SH[13]), .ZN(n505) );
  INV_X1 U367 ( .A(SH[31]), .ZN(n920) );
  AND2_X1 U368 ( .A1(n344), .A2(SH[1]), .ZN(n383) );
  NAND2_X1 U369 ( .A1(n241), .A2(SH[31]), .ZN(n344) );
  NAND4_X1 U370 ( .A1(n242), .A2(n244), .A3(n245), .A4(n243), .ZN(n241) );
  AND4_X1 U371 ( .A1(n249), .A2(SH[9]), .A3(SH[7]), .A4(SH[8]), .ZN(n242) );
  INV_X1 U372 ( .A(A[23]), .ZN(n952) );
  INV_X1 U374 ( .A(A[26]), .ZN(n949) );
  INV_X1 U375 ( .A(A[31]), .ZN(n944) );
  INV_X1 U376 ( .A(A[0]), .ZN(n974) );
  INV_X1 U377 ( .A(A[28]), .ZN(n947) );
  INV_X1 U378 ( .A(A[25]), .ZN(n950) );
  INV_X1 U379 ( .A(A[9]), .ZN(n966) );
  INV_X1 U380 ( .A(A[3]), .ZN(n972) );
  INV_X1 U381 ( .A(A[17]), .ZN(n958) );
  INV_X1 U382 ( .A(A[20]), .ZN(n955) );
  INV_X1 U383 ( .A(A[19]), .ZN(n956) );
  AND3_X1 U384 ( .A1(n248), .A2(SH[27]), .A3(n309), .ZN(n243) );
  AND2_X1 U385 ( .A1(SH[28]), .A2(SH[26]), .ZN(n309) );
  AND3_X1 U386 ( .A1(SH[24]), .A2(SH[23]), .A3(SH[25]), .ZN(n248) );
  INV_X1 U387 ( .A(A[16]), .ZN(n959) );
  NAND2_X1 U388 ( .A1(n915), .A2(A[30]), .ZN(n363) );
  INV_X1 U389 ( .A(A[24]), .ZN(n951) );
  NAND2_X1 U390 ( .A1(n939), .A2(A[29]), .ZN(n364) );
  INV_X1 U391 ( .A(A[13]), .ZN(n962) );
  INV_X1 U392 ( .A(A[22]), .ZN(n953) );
  INV_X1 U393 ( .A(A[12]), .ZN(n963) );
  NAND2_X1 U394 ( .A1(n935), .A2(A[15]), .ZN(n336) );
  INV_X1 U395 ( .A(A[27]), .ZN(n948) );
  AND3_X1 U396 ( .A1(SH[30]), .A2(SH[29]), .A3(SH[6]), .ZN(n249) );
  NAND2_X1 U397 ( .A1(n912), .A2(A[31]), .ZN(n362) );
  INV_X1 U398 ( .A(A[8]), .ZN(n967) );
  INV_X1 U399 ( .A(A[11]), .ZN(n964) );
  INV_X1 U400 ( .A(A[10]), .ZN(n965) );
  INV_X1 U401 ( .A(A[14]), .ZN(n961) );
  INV_X1 U402 ( .A(A[18]), .ZN(n957) );
  INV_X1 U403 ( .A(A[21]), .ZN(n954) );
  INV_X1 U404 ( .A(A[30]), .ZN(n945) );
  INV_X1 U405 ( .A(A[5]), .ZN(n970) );
  INV_X1 U406 ( .A(A[6]), .ZN(n969) );
  AND4_X1 U407 ( .A1(n247), .A2(SH[22]), .A3(SH[20]), .A4(SH[21]), .ZN(n244)
         );
  AND3_X1 U408 ( .A1(SH[18]), .A2(SH[17]), .A3(SH[19]), .ZN(n247) );
  INV_X1 U409 ( .A(A[4]), .ZN(n971) );
  INV_X1 U410 ( .A(A[7]), .ZN(n968) );
  OR3_X1 U411 ( .A1(SH[20]), .A2(SH[21]), .A3(SH[19]), .ZN(n257) );
  OR3_X1 U412 ( .A1(SH[14]), .A2(SH[15]), .A3(SH[13]), .ZN(n258) );
  OR2_X1 U413 ( .A1(n273), .A2(n960), .ZN(n358) );
  INV_X1 U414 ( .A(A[15]), .ZN(n960) );
  OR2_X1 U415 ( .A1(n946), .A2(n334), .ZN(n318) );
  INV_X1 U416 ( .A(A[29]), .ZN(n946) );
  OAI22_X1 U417 ( .A1(n189), .A2(n916), .B1(n190), .B2(n919), .ZN(B[16]) );
  OAI22_X1 U418 ( .A1(n125), .A2(n112), .B1(n126), .B2(n113), .ZN(B[29]) );
endmodule


module SHIFTER_M32_N5 ( A, B, LEFT_RIGHT, OUTPUT );
  input [31:0] A;
  input [31:0] B;
  output [31:0] OUTPUT;
  input LEFT_RIGHT;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298;

  SHIFTER_M32_N5_DW01_ash_0 sll_29 ( .A(A), .DATA_TC(1'b0), .SH(B), .SH_TC(
        1'b1), .B({N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, 
        N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37, N36, N35, N34}) );
  SHIFTER_M32_N5_DW_rash_0 srl_27 ( .A(A), .DATA_TC(1'b0), .SH(B), .SH_TC(1'b1), .B({N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
        N4, N3, N2}) );
  INV_X1 U1 ( .A(n298), .ZN(n288) );
  INV_X1 U2 ( .A(n298), .ZN(n289) );
  BUF_X1 U7 ( .A(n285), .Z(n290) );
  BUF_X1 U8 ( .A(n287), .Z(n297) );
  BUF_X1 U9 ( .A(n287), .Z(n296) );
  BUF_X1 U10 ( .A(n286), .Z(n295) );
  BUF_X1 U11 ( .A(n286), .Z(n294) );
  BUF_X1 U12 ( .A(n286), .Z(n293) );
  BUF_X1 U13 ( .A(n285), .Z(n292) );
  BUF_X1 U14 ( .A(n285), .Z(n291) );
  BUF_X1 U15 ( .A(n287), .Z(n298) );
  INV_X1 U16 ( .A(n46), .ZN(OUTPUT[5]) );
  AOI22_X1 U17 ( .A1(N7), .A2(n288), .B1(N39), .B2(n291), .ZN(n46) );
  INV_X1 U18 ( .A(n45), .ZN(OUTPUT[6]) );
  AOI22_X1 U19 ( .A1(N8), .A2(n289), .B1(N40), .B2(n290), .ZN(n45) );
  INV_X1 U20 ( .A(n44), .ZN(OUTPUT[7]) );
  AOI22_X1 U21 ( .A1(N9), .A2(n288), .B1(N41), .B2(n290), .ZN(n44) );
  INV_X1 U22 ( .A(n42), .ZN(OUTPUT[9]) );
  AOI22_X1 U23 ( .A1(N11), .A2(n289), .B1(N43), .B2(n290), .ZN(n42) );
  INV_X1 U24 ( .A(n49), .ZN(OUTPUT[31]) );
  AOI22_X1 U25 ( .A1(N33), .A2(n288), .B1(N65), .B2(n291), .ZN(n49) );
  INV_X1 U26 ( .A(n72), .ZN(OUTPUT[10]) );
  AOI22_X1 U27 ( .A1(N12), .A2(n288), .B1(N44), .B2(n297), .ZN(n72) );
  INV_X1 U28 ( .A(n58), .ZN(OUTPUT[23]) );
  AOI22_X1 U29 ( .A1(N25), .A2(n289), .B1(N57), .B2(n294), .ZN(n58) );
  INV_X1 U30 ( .A(n69), .ZN(OUTPUT[13]) );
  AOI22_X1 U31 ( .A1(N15), .A2(n288), .B1(N47), .B2(n296), .ZN(n69) );
  INV_X1 U32 ( .A(n70), .ZN(OUTPUT[12]) );
  AOI22_X1 U33 ( .A1(N14), .A2(n288), .B1(N46), .B2(n297), .ZN(n70) );
  INV_X1 U34 ( .A(n67), .ZN(OUTPUT[15]) );
  AOI22_X1 U35 ( .A1(N17), .A2(n288), .B1(N49), .B2(n296), .ZN(n67) );
  INV_X1 U36 ( .A(n65), .ZN(OUTPUT[17]) );
  AOI22_X1 U37 ( .A1(N19), .A2(n288), .B1(N51), .B2(n295), .ZN(n65) );
  INV_X1 U38 ( .A(n56), .ZN(OUTPUT[25]) );
  AOI22_X1 U39 ( .A1(N27), .A2(n289), .B1(N59), .B2(n293), .ZN(n56) );
  INV_X1 U40 ( .A(n55), .ZN(OUTPUT[26]) );
  AOI22_X1 U41 ( .A1(N28), .A2(n289), .B1(N60), .B2(n293), .ZN(n55) );
  INV_X1 U42 ( .A(n54), .ZN(OUTPUT[27]) );
  AOI22_X1 U43 ( .A1(N29), .A2(n289), .B1(N61), .B2(n293), .ZN(n54) );
  INV_X1 U44 ( .A(n71), .ZN(OUTPUT[11]) );
  AOI22_X1 U45 ( .A1(N13), .A2(n288), .B1(N45), .B2(n297), .ZN(n71) );
  INV_X1 U46 ( .A(n60), .ZN(OUTPUT[21]) );
  AOI22_X1 U47 ( .A1(N23), .A2(n289), .B1(N55), .B2(n294), .ZN(n60) );
  INV_X1 U48 ( .A(n62), .ZN(OUTPUT[1]) );
  AOI22_X1 U49 ( .A1(N3), .A2(n288), .B1(N35), .B2(n295), .ZN(n62) );
  INV_X1 U50 ( .A(n53), .ZN(OUTPUT[28]) );
  AOI22_X1 U51 ( .A1(N30), .A2(n289), .B1(N62), .B2(n292), .ZN(n53) );
  AOI22_X1 U52 ( .A1(N2), .A2(n288), .B1(N34), .B2(n297), .ZN(n73) );
  BUF_X1 U53 ( .A(LEFT_RIGHT), .Z(n287) );
  BUF_X1 U54 ( .A(LEFT_RIGHT), .Z(n286) );
  BUF_X1 U55 ( .A(LEFT_RIGHT), .Z(n285) );
  INV_X1 U56 ( .A(n48), .ZN(OUTPUT[3]) );
  AOI22_X1 U57 ( .A1(N5), .A2(n289), .B1(N37), .B2(n291), .ZN(n48) );
  INV_X1 U58 ( .A(n47), .ZN(OUTPUT[4]) );
  AOI22_X1 U59 ( .A1(N6), .A2(n288), .B1(N38), .B2(n291), .ZN(n47) );
  INV_X1 U60 ( .A(n43), .ZN(OUTPUT[8]) );
  AOI22_X1 U61 ( .A1(N10), .A2(n289), .B1(N42), .B2(n290), .ZN(n43) );
  INV_X1 U62 ( .A(n61), .ZN(OUTPUT[20]) );
  AOI22_X1 U63 ( .A1(N22), .A2(n289), .B1(N54), .B2(n294), .ZN(n61) );
  INV_X1 U64 ( .A(n68), .ZN(OUTPUT[14]) );
  AOI22_X1 U65 ( .A1(N16), .A2(n288), .B1(N48), .B2(n296), .ZN(n68) );
  INV_X1 U66 ( .A(n57), .ZN(OUTPUT[24]) );
  AOI22_X1 U67 ( .A1(N26), .A2(n289), .B1(N58), .B2(n293), .ZN(n57) );
  INV_X1 U68 ( .A(n59), .ZN(OUTPUT[22]) );
  AOI22_X1 U69 ( .A1(N24), .A2(n289), .B1(N56), .B2(n294), .ZN(n59) );
  INV_X1 U70 ( .A(n64), .ZN(OUTPUT[18]) );
  AOI22_X1 U71 ( .A1(N20), .A2(n288), .B1(N52), .B2(n295), .ZN(n64) );
  INV_X1 U72 ( .A(n63), .ZN(OUTPUT[19]) );
  AOI22_X1 U73 ( .A1(N21), .A2(n288), .B1(N53), .B2(n295), .ZN(n63) );
  INV_X1 U74 ( .A(n51), .ZN(OUTPUT[2]) );
  AOI22_X1 U75 ( .A1(N4), .A2(n289), .B1(N36), .B2(n292), .ZN(n51) );
  INV_X1 U76 ( .A(n50), .ZN(OUTPUT[30]) );
  AOI22_X1 U77 ( .A1(N32), .A2(n289), .B1(N64), .B2(n292), .ZN(n50) );
  INV_X1 U78 ( .A(n66), .ZN(OUTPUT[16]) );
  AOI22_X1 U79 ( .A1(N18), .A2(n288), .B1(N50), .B2(n296), .ZN(n66) );
  INV_X1 U80 ( .A(n52), .ZN(OUTPUT[29]) );
  AOI22_X1 U81 ( .A1(N31), .A2(n289), .B1(N63), .B2(n292), .ZN(n52) );
  INV_X1 U82 ( .A(n73), .ZN(OUTPUT[0]) );
endmodule


module PGnet_0 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_30 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_29 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_28 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_27 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_26 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_25 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_24 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_23 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_22 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_21 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_20 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_19 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_18 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_17 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_16 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_15 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_14 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_13 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_12 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_11 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_10 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_9 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_8 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_7 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_6 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_5 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_4 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_3 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_2 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_1 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module G_0 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n2;

  AOI21_X1 U1 ( .B1(p1), .B2(g2), .A(g1), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(g_Out) );
endmodule


module G_9 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module PG_0 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n2) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_26 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_25 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_24 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_23 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_22 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module PG_21 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module PG_20 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_19 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_18 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_17 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module PG_16 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_15 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_14 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module PG_13 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module G_8 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module PG_12 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module PG_11 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_10 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_9 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_8 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_7 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_6 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module G_7 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module PG_5 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_4 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module PG_3 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module G_6 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module G_5 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module PG_2 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module PG_1 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n16) );
endmodule


module G_4 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module G_3 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module G_2 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module G_1 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n16;

  INV_X1 U1 ( .A(n16), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n16) );
endmodule


module Cg ( A, B, cin0, cout );
  input [31:0] A;
  input [31:0] B;
  output [7:0] cout;
  input cin0;
  wire   n3, n6, n7, p0, g0, \gsignal[4][31] , \gsignal[4][27] ,
         \gsignal[3][31] , \gsignal[3][23] , \gsignal[3][15] ,
         \gsignal[2][31] , \gsignal[2][27] , \gsignal[2][23] ,
         \gsignal[2][19] , \gsignal[2][15] , \gsignal[2][11] , \gsignal[2][7] ,
         \gsignal[1][31] , \gsignal[1][29] , \gsignal[1][27] ,
         \gsignal[1][25] , \gsignal[1][23] , \gsignal[1][21] ,
         \gsignal[1][19] , \gsignal[1][17] , \gsignal[1][15] ,
         \gsignal[1][13] , \gsignal[1][11] , \gsignal[1][9] , \gsignal[1][7] ,
         \gsignal[1][5] , \gsignal[1][3] , \gsignal[1][1] , \gsignal[0][31] ,
         \gsignal[0][30] , \gsignal[0][29] , \gsignal[0][28] ,
         \gsignal[0][27] , \gsignal[0][26] , \gsignal[0][25] ,
         \gsignal[0][24] , \gsignal[0][23] , \gsignal[0][22] ,
         \gsignal[0][21] , \gsignal[0][20] , \gsignal[0][19] ,
         \gsignal[0][18] , \gsignal[0][17] , \gsignal[0][16] ,
         \gsignal[0][15] , \gsignal[0][14] , \gsignal[0][13] ,
         \gsignal[0][12] , \gsignal[0][11] , \gsignal[0][10] , \gsignal[0][9] ,
         \gsignal[0][8] , \gsignal[0][7] , \gsignal[0][6] , \gsignal[0][5] ,
         \gsignal[0][4] , \gsignal[0][3] , \gsignal[0][2] , \gsignal[0][1] ,
         \gsignal[0][0] , \psignal[4][31] , \psignal[4][27] , \psignal[3][31] ,
         \psignal[3][23] , \psignal[3][15] , \psignal[2][31] ,
         \psignal[2][27] , \psignal[2][23] , \psignal[2][19] ,
         \psignal[2][15] , \psignal[2][11] , \psignal[2][7] , \psignal[1][31] ,
         \psignal[1][29] , \psignal[1][27] , \psignal[1][25] ,
         \psignal[1][23] , \psignal[1][21] , \psignal[1][19] ,
         \psignal[1][17] , \psignal[1][15] , \psignal[1][13] ,
         \psignal[1][11] , \psignal[1][9] , \psignal[1][7] , \psignal[1][5] ,
         \psignal[1][3] , \psignal[0][31] , \psignal[0][30] , \psignal[0][29] ,
         \psignal[0][28] , \psignal[0][27] , \psignal[0][26] ,
         \psignal[0][25] , \psignal[0][24] , \psignal[0][23] ,
         \psignal[0][22] , \psignal[0][21] , \psignal[0][20] ,
         \psignal[0][19] , \psignal[0][18] , \psignal[0][17] ,
         \psignal[0][16] , \psignal[0][15] , \psignal[0][14] ,
         \psignal[0][13] , \psignal[0][12] , \psignal[0][11] ,
         \psignal[0][10] , \psignal[0][9] , \psignal[0][8] , \psignal[0][7] ,
         \psignal[0][6] , \psignal[0][5] , \psignal[0][4] , \psignal[0][3] ,
         \psignal[0][2] , \psignal[0][1] ;
  assign cout[3] = n3;
  assign cout[1] = n6;
  assign cout[0] = n7;

  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(p0) );
  PGnet_0 PGN1_31 ( .A(A[31]), .B(B[31]), .p(\psignal[0][31] ), .g(
        \gsignal[0][31] ) );
  PGnet_30 PGN1_30 ( .A(A[30]), .B(B[30]), .p(\psignal[0][30] ), .g(
        \gsignal[0][30] ) );
  PGnet_29 PGN1_29 ( .A(A[29]), .B(B[29]), .p(\psignal[0][29] ), .g(
        \gsignal[0][29] ) );
  PGnet_28 PGN1_28 ( .A(A[28]), .B(B[28]), .p(\psignal[0][28] ), .g(
        \gsignal[0][28] ) );
  PGnet_27 PGN1_27 ( .A(A[27]), .B(B[27]), .p(\psignal[0][27] ), .g(
        \gsignal[0][27] ) );
  PGnet_26 PGN1_26 ( .A(A[26]), .B(B[26]), .p(\psignal[0][26] ), .g(
        \gsignal[0][26] ) );
  PGnet_25 PGN1_25 ( .A(A[25]), .B(B[25]), .p(\psignal[0][25] ), .g(
        \gsignal[0][25] ) );
  PGnet_24 PGN1_24 ( .A(A[24]), .B(B[24]), .p(\psignal[0][24] ), .g(
        \gsignal[0][24] ) );
  PGnet_23 PGN1_23 ( .A(A[23]), .B(B[23]), .p(\psignal[0][23] ), .g(
        \gsignal[0][23] ) );
  PGnet_22 PGN1_22 ( .A(A[22]), .B(B[22]), .p(\psignal[0][22] ), .g(
        \gsignal[0][22] ) );
  PGnet_21 PGN1_21 ( .A(A[21]), .B(B[21]), .p(\psignal[0][21] ), .g(
        \gsignal[0][21] ) );
  PGnet_20 PGN1_20 ( .A(A[20]), .B(B[20]), .p(\psignal[0][20] ), .g(
        \gsignal[0][20] ) );
  PGnet_19 PGN1_19 ( .A(A[19]), .B(B[19]), .p(\psignal[0][19] ), .g(
        \gsignal[0][19] ) );
  PGnet_18 PGN1_18 ( .A(A[18]), .B(B[18]), .p(\psignal[0][18] ), .g(
        \gsignal[0][18] ) );
  PGnet_17 PGN1_17 ( .A(A[17]), .B(B[17]), .p(\psignal[0][17] ), .g(
        \gsignal[0][17] ) );
  PGnet_16 PGN1_16 ( .A(A[16]), .B(B[16]), .p(\psignal[0][16] ), .g(
        \gsignal[0][16] ) );
  PGnet_15 PGN1_15 ( .A(A[15]), .B(B[15]), .p(\psignal[0][15] ), .g(
        \gsignal[0][15] ) );
  PGnet_14 PGN1_14 ( .A(A[14]), .B(B[14]), .p(\psignal[0][14] ), .g(
        \gsignal[0][14] ) );
  PGnet_13 PGN1_13 ( .A(A[13]), .B(B[13]), .p(\psignal[0][13] ), .g(
        \gsignal[0][13] ) );
  PGnet_12 PGN1_12 ( .A(A[12]), .B(B[12]), .p(\psignal[0][12] ), .g(
        \gsignal[0][12] ) );
  PGnet_11 PGN1_11 ( .A(A[11]), .B(B[11]), .p(\psignal[0][11] ), .g(
        \gsignal[0][11] ) );
  PGnet_10 PGN1_10 ( .A(A[10]), .B(B[10]), .p(\psignal[0][10] ), .g(
        \gsignal[0][10] ) );
  PGnet_9 PGN1_9 ( .A(A[9]), .B(B[9]), .p(\psignal[0][9] ), .g(\gsignal[0][9] ) );
  PGnet_8 PGN1_8 ( .A(A[8]), .B(B[8]), .p(\psignal[0][8] ), .g(\gsignal[0][8] ) );
  PGnet_7 PGN1_7 ( .A(A[7]), .B(B[7]), .p(\psignal[0][7] ), .g(\gsignal[0][7] ) );
  PGnet_6 PGN1_6 ( .A(A[6]), .B(B[6]), .p(\psignal[0][6] ), .g(\gsignal[0][6] ) );
  PGnet_5 PGN1_5 ( .A(A[5]), .B(B[5]), .p(\psignal[0][5] ), .g(\gsignal[0][5] ) );
  PGnet_4 PGN1_4 ( .A(A[4]), .B(B[4]), .p(\psignal[0][4] ), .g(\gsignal[0][4] ) );
  PGnet_3 PGN1_3 ( .A(A[3]), .B(B[3]), .p(\psignal[0][3] ), .g(\gsignal[0][3] ) );
  PGnet_2 PGN1_2 ( .A(A[2]), .B(B[2]), .p(\psignal[0][2] ), .g(\gsignal[0][2] ) );
  PGnet_1 PGN1_1 ( .A(A[1]), .B(B[1]), .p(\psignal[0][1] ), .g(\gsignal[0][1] ) );
  G_0 PGN0_0 ( .p1(p0), .g1(g0), .g2(cin0), .g_Out(\gsignal[0][0] ) );
  G_9 g0_0_1 ( .p1(\psignal[0][1] ), .g1(\gsignal[0][1] ), .g2(\gsignal[0][0] ), .g_Out(\gsignal[1][1] ) );
  PG_0 PGelements_0_3 ( .p1(\psignal[0][3] ), .g1(\gsignal[0][3] ), .p2(
        \psignal[0][2] ), .g2(\gsignal[0][2] ), .p_Out(\psignal[1][3] ), 
        .g_Out(\gsignal[1][3] ) );
  PG_26 PGelements_0_5 ( .p1(\psignal[0][5] ), .g1(\gsignal[0][5] ), .p2(
        \psignal[0][4] ), .g2(\gsignal[0][4] ), .p_Out(\psignal[1][5] ), 
        .g_Out(\gsignal[1][5] ) );
  PG_25 PGelements_0_7 ( .p1(\psignal[0][7] ), .g1(\gsignal[0][7] ), .p2(
        \psignal[0][6] ), .g2(\gsignal[0][6] ), .p_Out(\psignal[1][7] ), 
        .g_Out(\gsignal[1][7] ) );
  PG_24 PGelements_0_9 ( .p1(\psignal[0][9] ), .g1(\gsignal[0][9] ), .p2(
        \psignal[0][8] ), .g2(\gsignal[0][8] ), .p_Out(\psignal[1][9] ), 
        .g_Out(\gsignal[1][9] ) );
  PG_23 PGelements_0_11 ( .p1(\psignal[0][11] ), .g1(\gsignal[0][11] ), .p2(
        \psignal[0][10] ), .g2(\gsignal[0][10] ), .p_Out(\psignal[1][11] ), 
        .g_Out(\gsignal[1][11] ) );
  PG_22 PGelements_0_13 ( .p1(\psignal[0][13] ), .g1(\gsignal[0][13] ), .p2(
        \psignal[0][12] ), .g2(\gsignal[0][12] ), .p_Out(\psignal[1][13] ), 
        .g_Out(\gsignal[1][13] ) );
  PG_21 PGelements_0_15 ( .p1(\psignal[0][15] ), .g1(\gsignal[0][15] ), .p2(
        \psignal[0][14] ), .g2(\gsignal[0][14] ), .p_Out(\psignal[1][15] ), 
        .g_Out(\gsignal[1][15] ) );
  PG_20 PGelements_0_17 ( .p1(\psignal[0][17] ), .g1(\gsignal[0][17] ), .p2(
        \psignal[0][16] ), .g2(\gsignal[0][16] ), .p_Out(\psignal[1][17] ), 
        .g_Out(\gsignal[1][17] ) );
  PG_19 PGelements_0_19 ( .p1(\psignal[0][19] ), .g1(\gsignal[0][19] ), .p2(
        \psignal[0][18] ), .g2(\gsignal[0][18] ), .p_Out(\psignal[1][19] ), 
        .g_Out(\gsignal[1][19] ) );
  PG_18 PGelements_0_21 ( .p1(\psignal[0][21] ), .g1(\gsignal[0][21] ), .p2(
        \psignal[0][20] ), .g2(\gsignal[0][20] ), .p_Out(\psignal[1][21] ), 
        .g_Out(\gsignal[1][21] ) );
  PG_17 PGelements_0_23 ( .p1(\psignal[0][23] ), .g1(\gsignal[0][23] ), .p2(
        \psignal[0][22] ), .g2(\gsignal[0][22] ), .p_Out(\psignal[1][23] ), 
        .g_Out(\gsignal[1][23] ) );
  PG_16 PGelements_0_25 ( .p1(\psignal[0][25] ), .g1(\gsignal[0][25] ), .p2(
        \psignal[0][24] ), .g2(\gsignal[0][24] ), .p_Out(\psignal[1][25] ), 
        .g_Out(\gsignal[1][25] ) );
  PG_15 PGelements_0_27 ( .p1(\psignal[0][27] ), .g1(\gsignal[0][27] ), .p2(
        \psignal[0][26] ), .g2(\gsignal[0][26] ), .p_Out(\psignal[1][27] ), 
        .g_Out(\gsignal[1][27] ) );
  PG_14 PGelements_0_29 ( .p1(\psignal[0][29] ), .g1(\gsignal[0][29] ), .p2(
        \psignal[0][28] ), .g2(\gsignal[0][28] ), .p_Out(\psignal[1][29] ), 
        .g_Out(\gsignal[1][29] ) );
  PG_13 PGelements_0_31 ( .p1(\psignal[0][31] ), .g1(\gsignal[0][31] ), .p2(
        \psignal[0][30] ), .g2(\gsignal[0][30] ), .p_Out(\psignal[1][31] ), 
        .g_Out(\gsignal[1][31] ) );
  G_8 g0_1_3 ( .p1(\psignal[1][3] ), .g1(\gsignal[1][3] ), .g2(\gsignal[1][1] ), .g_Out(n7) );
  PG_12 PGelements_1_7 ( .p1(\psignal[1][7] ), .g1(\gsignal[1][7] ), .p2(
        \psignal[1][5] ), .g2(\gsignal[1][5] ), .p_Out(\psignal[2][7] ), 
        .g_Out(\gsignal[2][7] ) );
  PG_11 PGelements_1_11 ( .p1(\psignal[1][11] ), .g1(\gsignal[1][11] ), .p2(
        \psignal[1][9] ), .g2(\gsignal[1][9] ), .p_Out(\psignal[2][11] ), 
        .g_Out(\gsignal[2][11] ) );
  PG_10 PGelements_1_15 ( .p1(\psignal[1][15] ), .g1(\gsignal[1][15] ), .p2(
        \psignal[1][13] ), .g2(\gsignal[1][13] ), .p_Out(\psignal[2][15] ), 
        .g_Out(\gsignal[2][15] ) );
  PG_9 PGelements_1_19 ( .p1(\psignal[1][19] ), .g1(\gsignal[1][19] ), .p2(
        \psignal[1][17] ), .g2(\gsignal[1][17] ), .p_Out(\psignal[2][19] ), 
        .g_Out(\gsignal[2][19] ) );
  PG_8 PGelements_1_23 ( .p1(\psignal[1][23] ), .g1(\gsignal[1][23] ), .p2(
        \psignal[1][21] ), .g2(\gsignal[1][21] ), .p_Out(\psignal[2][23] ), 
        .g_Out(\gsignal[2][23] ) );
  PG_7 PGelements_1_27 ( .p1(\psignal[1][27] ), .g1(\gsignal[1][27] ), .p2(
        \psignal[1][25] ), .g2(\gsignal[1][25] ), .p_Out(\psignal[2][27] ), 
        .g_Out(\gsignal[2][27] ) );
  PG_6 PGelements_1_31 ( .p1(\psignal[1][31] ), .g1(\gsignal[1][31] ), .p2(
        \psignal[1][29] ), .g2(\gsignal[1][29] ), .p_Out(\psignal[2][31] ), 
        .g_Out(\gsignal[2][31] ) );
  G_7 g0_2_7 ( .p1(\psignal[2][7] ), .g1(\gsignal[2][7] ), .g2(n7), .g_Out(n6)
         );
  PG_5 PGelements_2_15 ( .p1(\psignal[2][15] ), .g1(\gsignal[2][15] ), .p2(
        \psignal[2][11] ), .g2(\gsignal[2][11] ), .p_Out(\psignal[3][15] ), 
        .g_Out(\gsignal[3][15] ) );
  PG_4 PGelements_2_23 ( .p1(\psignal[2][23] ), .g1(\gsignal[2][23] ), .p2(
        \psignal[2][19] ), .g2(\gsignal[2][19] ), .p_Out(\psignal[3][23] ), 
        .g_Out(\gsignal[3][23] ) );
  PG_3 PGelements_2_31 ( .p1(\psignal[2][31] ), .g1(\gsignal[2][31] ), .p2(
        \psignal[2][27] ), .g2(\gsignal[2][27] ), .p_Out(\psignal[3][31] ), 
        .g_Out(\gsignal[3][31] ) );
  G_6 g1_3_11 ( .p1(\psignal[2][11] ), .g1(\gsignal[2][11] ), .g2(n6), .g_Out(
        cout[2]) );
  G_5 g1_3_15 ( .p1(\psignal[3][15] ), .g1(\gsignal[3][15] ), .g2(n6), .g_Out(
        n3) );
  PG_2 pg1_3_27 ( .p1(\psignal[2][27] ), .g1(\gsignal[2][27] ), .p2(
        \psignal[3][15] ), .g2(\gsignal[3][15] ), .p_Out(\psignal[4][27] ), 
        .g_Out(\gsignal[4][27] ) );
  PG_1 pg1_3_31 ( .p1(\psignal[3][31] ), .g1(\gsignal[3][31] ), .p2(
        \psignal[3][15] ), .g2(\gsignal[3][15] ), .p_Out(\psignal[4][31] ), 
        .g_Out(\gsignal[4][31] ) );
  G_4 g1_4_19 ( .p1(\psignal[2][19] ), .g1(\gsignal[2][19] ), .g2(n3), .g_Out(
        cout[4]) );
  G_3 g1_4_23 ( .p1(\psignal[3][23] ), .g1(\gsignal[3][23] ), .g2(n3), .g_Out(
        cout[5]) );
  G_2 g1_4_27 ( .p1(\psignal[4][27] ), .g1(\gsignal[4][27] ), .g2(n3), .g_Out(
        cout[6]) );
  G_1 g1_4_31 ( .p1(\psignal[4][31] ), .g1(\gsignal[4][31] ), .g2(n3), .g_Out(
        cout[7]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(g0) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n2) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_6 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n6, n7, n8, n9, n52;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(ci), .ZN(n52) );
  INV_X1 U4 ( .A(n7), .ZN(s[2]) );
  AOI22_X1 U5 ( .A1(out0[2]), .A2(n52), .B1(out1[2]), .B2(ci), .ZN(n7) );
  INV_X1 U6 ( .A(n6), .ZN(s[3]) );
  AOI22_X1 U7 ( .A1(out0[3]), .A2(n52), .B1(out1[3]), .B2(ci), .ZN(n6) );
  INV_X1 U8 ( .A(n8), .ZN(s[1]) );
  AOI22_X1 U9 ( .A1(out0[1]), .A2(n52), .B1(out1[1]), .B2(ci), .ZN(n8) );
  INV_X1 U10 ( .A(n9), .ZN(s[0]) );
  AOI22_X1 U11 ( .A1(out0[0]), .A2(n52), .B1(out1[0]), .B2(ci), .ZN(n9) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_5 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n6, n7, n8, n9, n52;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(ci), .ZN(n52) );
  INV_X1 U4 ( .A(n6), .ZN(s[3]) );
  AOI22_X1 U5 ( .A1(out0[3]), .A2(n52), .B1(out1[3]), .B2(ci), .ZN(n6) );
  INV_X1 U6 ( .A(n7), .ZN(s[2]) );
  AOI22_X1 U7 ( .A1(out0[2]), .A2(n52), .B1(out1[2]), .B2(ci), .ZN(n7) );
  INV_X1 U8 ( .A(n8), .ZN(s[1]) );
  AOI22_X1 U9 ( .A1(out0[1]), .A2(n52), .B1(out1[1]), .B2(ci), .ZN(n8) );
  INV_X1 U10 ( .A(n9), .ZN(s[0]) );
  AOI22_X1 U11 ( .A1(out0[0]), .A2(n52), .B1(out1[0]), .B2(ci), .ZN(n9) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_4 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n52, n53, n54, n55, n56;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(ci), .ZN(n52) );
  INV_X1 U4 ( .A(n55), .ZN(s[2]) );
  AOI22_X1 U5 ( .A1(out0[2]), .A2(n52), .B1(out1[2]), .B2(ci), .ZN(n55) );
  INV_X1 U6 ( .A(n56), .ZN(s[3]) );
  AOI22_X1 U7 ( .A1(out0[3]), .A2(n52), .B1(out1[3]), .B2(ci), .ZN(n56) );
  INV_X1 U8 ( .A(n54), .ZN(s[1]) );
  AOI22_X1 U9 ( .A1(out0[1]), .A2(n52), .B1(out1[1]), .B2(ci), .ZN(n54) );
  INV_X1 U10 ( .A(n53), .ZN(s[0]) );
  AOI22_X1 U11 ( .A1(out0[0]), .A2(n52), .B1(out1[0]), .B2(ci), .ZN(n53) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_3 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n52, n53, n54, n55, n56;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(ci), .ZN(n52) );
  INV_X1 U4 ( .A(n55), .ZN(s[2]) );
  AOI22_X1 U5 ( .A1(out0[2]), .A2(n52), .B1(out1[2]), .B2(ci), .ZN(n55) );
  INV_X1 U6 ( .A(n56), .ZN(s[3]) );
  AOI22_X1 U7 ( .A1(out0[3]), .A2(n52), .B1(out1[3]), .B2(ci), .ZN(n56) );
  INV_X1 U8 ( .A(n54), .ZN(s[1]) );
  AOI22_X1 U9 ( .A1(out0[1]), .A2(n52), .B1(out1[1]), .B2(ci), .ZN(n54) );
  INV_X1 U10 ( .A(n53), .ZN(s[0]) );
  AOI22_X1 U11 ( .A1(out0[0]), .A2(n52), .B1(out1[0]), .B2(ci), .ZN(n53) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_2 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n52, n53, n54, n55, n56;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(ci), .ZN(n52) );
  INV_X1 U4 ( .A(n55), .ZN(s[2]) );
  AOI22_X1 U5 ( .A1(out0[2]), .A2(n52), .B1(out1[2]), .B2(ci), .ZN(n55) );
  INV_X1 U6 ( .A(n56), .ZN(s[3]) );
  AOI22_X1 U7 ( .A1(out0[3]), .A2(n52), .B1(out1[3]), .B2(ci), .ZN(n56) );
  INV_X1 U8 ( .A(n54), .ZN(s[1]) );
  AOI22_X1 U9 ( .A1(out0[1]), .A2(n52), .B1(out1[1]), .B2(ci), .ZN(n54) );
  INV_X1 U10 ( .A(n53), .ZN(s[0]) );
  AOI22_X1 U11 ( .A1(out0[0]), .A2(n52), .B1(out1[0]), .B2(ci), .ZN(n53) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n23, n24;

  XOR2_X1 U3 ( .A(Ci), .B(n23), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n23) );
  INV_X1 U1 ( .A(n24), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n23), .B2(Ci), .ZN(n24) );
endmodule


module RCA_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_1 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n52, n53, n54, n55, n56;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(ci), .ZN(n52) );
  INV_X1 U4 ( .A(n55), .ZN(s[2]) );
  AOI22_X1 U5 ( .A1(out0[2]), .A2(n52), .B1(out1[2]), .B2(ci), .ZN(n55) );
  INV_X1 U6 ( .A(n56), .ZN(s[3]) );
  AOI22_X1 U7 ( .A1(out0[3]), .A2(n52), .B1(out1[3]), .B2(ci), .ZN(n56) );
  INV_X1 U8 ( .A(n54), .ZN(s[1]) );
  AOI22_X1 U9 ( .A1(out0[1]), .A2(n52), .B1(out1[1]), .B2(ci), .ZN(n54) );
  INV_X1 U10 ( .A(n53), .ZN(s[0]) );
  AOI22_X1 U11 ( .A1(out0[0]), .A2(n52), .B1(out1[0]), .B2(ci), .ZN(n53) );
endmodule


module CSA ( A, B, c, s );
  input [31:0] A;
  input [31:0] B;
  input [7:0] c;
  output [31:0] s;


  CSb_0 CSbi_0 ( .A(A[3:0]), .B(B[3:0]), .ci(c[0]), .s(s[3:0]) );
  CSb_7 CSbi_1 ( .A(A[7:4]), .B(B[7:4]), .ci(c[1]), .s(s[7:4]) );
  CSb_6 CSbi_2 ( .A(A[11:8]), .B(B[11:8]), .ci(c[2]), .s(s[11:8]) );
  CSb_5 CSbi_3 ( .A(A[15:12]), .B(B[15:12]), .ci(c[3]), .s(s[15:12]) );
  CSb_4 CSbi_4 ( .A(A[19:16]), .B(B[19:16]), .ci(c[4]), .s(s[19:16]) );
  CSb_3 CSbi_5 ( .A(A[23:20]), .B(B[23:20]), .ci(c[5]), .s(s[23:20]) );
  CSb_2 CSbi_6 ( .A(A[27:24]), .B(B[27:24]), .ci(c[6]), .s(s[27:24]) );
  CSb_1 CSbi_7 ( .A(A[31:28]), .B(B[31:28]), .ci(c[7]), .s(s[31:28]) );
endmodule


module P4ADDER_n_bit32 ( A, B, cin0, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input cin0;
  wire   n1, n5, n6, n7, n20, n21;
  wire   [7:1] carries;
  wire   [31:0] BS;
  wire   SYNOPSYS_UNCONNECTED__0;

  XOR2_X1 U1 ( .A(n21), .B(B[13]), .Z(n7) );
  XOR2_X1 U2 ( .A(n21), .B(B[7]), .Z(n6) );
  XOR2_X1 U3 ( .A(n21), .B(B[14]), .Z(n5) );
  XOR2_X1 U4 ( .A(n21), .B(B[0]), .Z(n1) );
  XOR2_X1 U5 ( .A(n21), .B(B[9]), .Z(BS[9]) );
  XOR2_X1 U6 ( .A(n21), .B(B[8]), .Z(BS[8]) );
  XOR2_X1 U7 ( .A(n21), .B(B[6]), .Z(BS[6]) );
  XOR2_X1 U8 ( .A(n21), .B(B[5]), .Z(BS[5]) );
  XOR2_X1 U9 ( .A(n21), .B(B[4]), .Z(BS[4]) );
  XOR2_X1 U10 ( .A(n21), .B(B[3]), .Z(BS[3]) );
  XOR2_X1 U11 ( .A(n21), .B(B[31]), .Z(BS[31]) );
  XOR2_X1 U12 ( .A(n21), .B(B[30]), .Z(BS[30]) );
  XOR2_X1 U13 ( .A(n21), .B(B[2]), .Z(BS[2]) );
  XOR2_X1 U14 ( .A(n21), .B(B[29]), .Z(BS[29]) );
  XOR2_X1 U15 ( .A(n21), .B(B[28]), .Z(BS[28]) );
  XOR2_X1 U16 ( .A(n20), .B(B[27]), .Z(BS[27]) );
  XOR2_X1 U17 ( .A(n20), .B(B[26]), .Z(BS[26]) );
  XOR2_X1 U18 ( .A(n20), .B(B[25]), .Z(BS[25]) );
  XOR2_X1 U19 ( .A(n20), .B(B[24]), .Z(BS[24]) );
  XOR2_X1 U20 ( .A(n20), .B(B[23]), .Z(BS[23]) );
  XOR2_X1 U21 ( .A(n20), .B(B[22]), .Z(BS[22]) );
  XOR2_X1 U22 ( .A(n20), .B(B[21]), .Z(BS[21]) );
  XOR2_X1 U23 ( .A(n20), .B(B[20]), .Z(BS[20]) );
  XOR2_X1 U24 ( .A(n20), .B(B[1]), .Z(BS[1]) );
  XOR2_X1 U25 ( .A(n20), .B(B[19]), .Z(BS[19]) );
  XOR2_X1 U26 ( .A(n20), .B(B[18]), .Z(BS[18]) );
  XOR2_X1 U27 ( .A(n20), .B(B[17]), .Z(BS[17]) );
  XOR2_X1 U28 ( .A(n20), .B(B[16]), .Z(BS[16]) );
  XOR2_X1 U29 ( .A(n20), .B(B[15]), .Z(BS[15]) );
  XOR2_X1 U30 ( .A(n20), .B(B[12]), .Z(BS[12]) );
  XOR2_X1 U31 ( .A(n20), .B(B[11]), .Z(BS[11]) );
  XOR2_X1 U32 ( .A(n21), .B(B[10]), .Z(BS[10]) );
  Cg CG1 ( .A(A), .B({BS[31:15], n5, n7, BS[12:8], n6, BS[6:1], n1}), .cin0(
        n20), .cout({SYNOPSYS_UNCONNECTED__0, carries}) );
  CSA CSA1 ( .A(A), .B({BS[31:15], n5, n7, BS[12:8], n6, BS[6:1], n1}), .c({
        carries, n21}), .s(S) );
  BUF_X1 U33 ( .A(cin0), .Z(n20) );
  BUF_X1 U34 ( .A(cin0), .Z(n21) );
endmodule


module COMPARATOR_M32_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n26, n27, n29, n30, n31, n32, n33, n34,
         n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n55, n56, n58, n59, n60, n61, n62, n63, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n82, n83,
         n86, n88, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n100,
         n101, n103, n105, n106, n107, n108, n109, n110, n111, n112, n115,
         n116, n118, n119, n120, n121, n122, n123, n124, n125, n126, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n141,
         n142, n144, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n159, n161, n162, n163, n164, n165, n167, n168, n169,
         n172, n175, n176, n177, n178, n179, n180, n181, n182, n183, n193,
         n194, n195, n198, n200, n201, n204, n206, n207, n208, n209, n210,
         n211, n212, n216, n218, n225, n226, n227, n228, n231, n233, n234,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n255, n256,
         n257, n258, n263, n264, n268, n269, n270, n271, n272, n273, n276,
         n278, n286, n287, n288, n289, n290, n292, n293, n294, n295, n298,
         n300, n301, n303, n305, n306, n313, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907;

  NAND3_X1 U281 ( .A1(n16), .A2(n17), .A3(n15), .ZN(n11) );
  NAND3_X1 U282 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n20) );
  NAND3_X1 U283 ( .A1(n818), .A2(n29), .A3(n813), .ZN(n22) );
  NAND3_X1 U284 ( .A1(n39), .A2(n826), .A3(n40), .ZN(n43) );
  NAND3_X1 U285 ( .A1(n40), .A2(n52), .A3(n53), .ZN(n51) );
  NAND3_X1 U286 ( .A1(n831), .A2(n58), .A3(n827), .ZN(n52) );
  NAND3_X1 U287 ( .A1(n60), .A2(n39), .A3(n61), .ZN(n50) );
  NAND3_X1 U288 ( .A1(n76), .A2(n77), .A3(n78), .ZN(n75) );
  NAND3_X1 U289 ( .A1(n97), .A2(n854), .A3(n98), .ZN(n101) );
  NAND3_X1 U292 ( .A1(n859), .A2(n855), .A3(n118), .ZN(n111) );
  NAND3_X1 U293 ( .A1(n120), .A2(n97), .A3(n121), .ZN(n109) );
  NAND3_X1 U294 ( .A1(n132), .A2(n137), .A3(n138), .ZN(n123) );
  NAND3_X1 U295 ( .A1(n872), .A2(n144), .A3(n868), .ZN(n137) );
  NAND3_X1 U296 ( .A1(n151), .A2(n152), .A3(n153), .ZN(n147) );
  NAND3_X1 U297 ( .A1(n167), .A2(n168), .A3(n169), .ZN(n164) );
  NAND3_X1 U298 ( .A1(n27), .A2(n813), .A3(n820), .ZN(n167) );
  NAND3_X1 U299 ( .A1(n183), .A2(n824), .A3(n46), .ZN(n182) );
  NAND3_X1 U300 ( .A1(n183), .A2(n46), .A3(n41), .ZN(n180) );
  NAND3_X1 U301 ( .A1(n833), .A2(n56), .A3(n827), .ZN(n195) );
  NAND3_X1 U304 ( .A1(n216), .A2(n70), .A3(n72), .ZN(n211) );
  NAND3_X1 U305 ( .A1(n218), .A2(n1), .A3(n827), .ZN(n209) );
  NAND3_X1 U307 ( .A1(n216), .A2(n838), .A3(n70), .ZN(n218) );
  NAND3_X1 U308 ( .A1(n245), .A2(n852), .A3(n105), .ZN(n244) );
  NAND3_X1 U309 ( .A1(n245), .A2(n105), .A3(n99), .ZN(n242) );
  NAND3_X1 U310 ( .A1(n862), .A2(n116), .A3(n855), .ZN(n257) );
  NAND3_X1 U311 ( .A1(n276), .A2(n136), .A3(n133), .ZN(n272) );
  NAND3_X1 U312 ( .A1(n278), .A2(n860), .A3(n855), .ZN(n270) );
  NAND3_X1 U313 ( .A1(n276), .A2(n866), .A3(n136), .ZN(n278) );
  NAND3_X1 U314 ( .A1(n286), .A2(n287), .A3(n288), .ZN(n268) );
  NAND3_X1 U315 ( .A1(n293), .A2(n294), .A3(n295), .ZN(n287) );
  AOI21_X1 U1 ( .B1(n238), .B2(n239), .A(n240), .ZN(n206) );
  NAND2_X1 U2 ( .A1(n268), .A2(n269), .ZN(n238) );
  NOR2_X1 U3 ( .A1(n255), .A2(n256), .ZN(n239) );
  NAND4_X1 U4 ( .A1(n241), .A2(n242), .A3(n243), .A4(n244), .ZN(n240) );
  AOI21_X1 U5 ( .B1(n176), .B2(n177), .A(n178), .ZN(n163) );
  AND3_X1 U6 ( .A1(n193), .A2(n194), .A3(n195), .ZN(n177) );
  NAND4_X1 U7 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(n178) );
  OAI21_X1 U8 ( .B1(n206), .B2(n207), .A(n208), .ZN(n176) );
  OAI21_X1 U9 ( .B1(n47), .B2(n48), .A(n49), .ZN(n18) );
  NAND2_X1 U10 ( .A1(n62), .A2(n63), .ZN(n48) );
  NOR2_X1 U11 ( .A1(n50), .A2(n51), .ZN(n49) );
  AOI21_X1 U12 ( .B1(n73), .B2(n74), .A(n75), .ZN(n47) );
  INV_X1 U13 ( .A(n55), .ZN(n827) );
  NOR2_X1 U14 ( .A1(n96), .A2(n83), .ZN(n243) );
  NOR2_X1 U15 ( .A1(n38), .A2(n26), .ZN(n181) );
  NOR2_X1 U16 ( .A1(n91), .A2(n92), .ZN(n74) );
  NAND2_X1 U17 ( .A1(n100), .A2(n101), .ZN(n91) );
  OAI21_X1 U18 ( .B1(n850), .B2(n94), .A(n95), .ZN(n92) );
  NOR2_X1 U19 ( .A1(n845), .A2(n849), .ZN(n100) );
  NOR2_X1 U20 ( .A1(n834), .A2(n829), .ZN(n212) );
  NOR2_X1 U21 ( .A1(n83), .A2(n845), .ZN(n79) );
  INV_X1 U22 ( .A(n26), .ZN(n813) );
  NOR2_X1 U23 ( .A1(n96), .A2(n83), .ZN(n95) );
  NOR2_X1 U24 ( .A1(n38), .A2(n26), .ZN(n37) );
  NOR2_X1 U25 ( .A1(n130), .A2(n115), .ZN(n129) );
  NAND2_X1 U26 ( .A1(n843), .A2(n841), .ZN(n77) );
  NOR2_X1 U27 ( .A1(n840), .A2(n88), .ZN(n76) );
  AOI21_X1 U28 ( .B1(n79), .B2(n846), .A(n834), .ZN(n78) );
  INV_X1 U29 ( .A(n115), .ZN(n855) );
  NOR2_X1 U30 ( .A1(n141), .A2(n154), .ZN(n153) );
  NOR2_X1 U31 ( .A1(n141), .A2(n154), .ZN(n295) );
  INV_X1 U32 ( .A(n83), .ZN(n841) );
  INV_X1 U33 ( .A(n141), .ZN(n868) );
  NAND2_X1 U34 ( .A1(n107), .A2(n108), .ZN(n73) );
  NOR2_X1 U35 ( .A1(n109), .A2(n110), .ZN(n108) );
  OAI21_X1 U36 ( .B1(n122), .B2(n123), .A(n124), .ZN(n107) );
  NAND2_X1 U37 ( .A1(n111), .A2(n112), .ZN(n110) );
  INV_X1 U38 ( .A(n8), .ZN(LE) );
  INV_X1 U39 ( .A(n41), .ZN(n822) );
  INV_X1 U40 ( .A(n99), .ZN(n850) );
  INV_X1 U41 ( .A(n130), .ZN(n860) );
  NOR2_X1 U42 ( .A1(n9), .A2(n8), .ZN(EQ) );
  OAI21_X1 U43 ( .B1(n10), .B2(n11), .A(n12), .ZN(n8) );
  NOR2_X1 U44 ( .A1(n13), .A2(n3), .ZN(n12) );
  AOI21_X1 U45 ( .B1(n18), .B2(n19), .A(n20), .ZN(n10) );
  NAND2_X1 U46 ( .A1(n90), .A2(n231), .ZN(n83) );
  NAND2_X1 U47 ( .A1(n150), .A2(n298), .ZN(n141) );
  NAND2_X1 U48 ( .A1(n32), .A2(n172), .ZN(n26) );
  INV_X1 U49 ( .A(n45), .ZN(n826) );
  INV_X1 U50 ( .A(n103), .ZN(n854) );
  INV_X1 U51 ( .A(n120), .ZN(n852) );
  INV_X1 U52 ( .A(n60), .ZN(n824) );
  NAND4_X1 U53 ( .A1(n105), .A2(n103), .A3(n245), .A4(n264), .ZN(n255) );
  NOR2_X1 U54 ( .A1(n270), .A2(n271), .ZN(n269) );
  NAND2_X1 U55 ( .A1(n272), .A2(n273), .ZN(n271) );
  AND2_X1 U56 ( .A1(n132), .A2(n116), .ZN(n273) );
  NOR2_X1 U57 ( .A1(n33), .A2(n34), .ZN(n19) );
  NAND2_X1 U58 ( .A1(n42), .A2(n43), .ZN(n33) );
  OAI21_X1 U59 ( .B1(n822), .B2(n36), .A(n37), .ZN(n34) );
  AND2_X1 U60 ( .A1(n29), .A2(n46), .ZN(n42) );
  NAND2_X1 U61 ( .A1(n121), .A2(n264), .ZN(n115) );
  NOR2_X1 U62 ( .A1(n83), .A2(n106), .ZN(n234) );
  NOR2_X1 U63 ( .A1(n141), .A2(n144), .ZN(n290) );
  NOR2_X1 U64 ( .A1(n836), .A2(n65), .ZN(n63) );
  INV_X1 U65 ( .A(n70), .ZN(n836) );
  OAI21_X1 U66 ( .B1(n66), .B2(n67), .A(n58), .ZN(n65) );
  NAND2_X1 U67 ( .A1(n68), .A2(n69), .ZN(n67) );
  NOR2_X1 U68 ( .A1(n141), .A2(n292), .ZN(n289) );
  NAND2_X1 U69 ( .A1(n829), .A2(n827), .ZN(n53) );
  INV_X1 U70 ( .A(n59), .ZN(n831) );
  NAND2_X1 U71 ( .A1(n870), .A2(n868), .ZN(n138) );
  INV_X1 U72 ( .A(n142), .ZN(n870) );
  AND2_X1 U73 ( .A1(n16), .A2(n172), .ZN(n168) );
  NAND2_X1 U74 ( .A1(n817), .A2(n813), .ZN(n169) );
  NOR2_X1 U75 ( .A1(n209), .A2(n210), .ZN(n208) );
  NAND2_X1 U76 ( .A1(n211), .A2(n212), .ZN(n210) );
  NOR2_X1 U77 ( .A1(n125), .A2(n126), .ZN(n124) );
  OAI21_X1 U78 ( .B1(n864), .B2(n128), .A(n129), .ZN(n126) );
  OAI211_X1 U79 ( .C1(n134), .C2(n135), .A(n118), .B(n136), .ZN(n125) );
  INV_X1 U80 ( .A(n133), .ZN(n864) );
  NOR2_X1 U81 ( .A1(n843), .A2(n237), .ZN(n233) );
  AND2_X1 U82 ( .A1(n31), .A2(n32), .ZN(n21) );
  NAND2_X1 U83 ( .A1(n815), .A2(n813), .ZN(n23) );
  INV_X1 U84 ( .A(n119), .ZN(n859) );
  NOR2_X1 U85 ( .A1(n2), .A2(n71), .ZN(n62) );
  NAND2_X1 U86 ( .A1(n827), .A2(n1), .ZN(n71) );
  AND3_X1 U87 ( .A1(n69), .A2(n68), .A3(n72), .ZN(n2) );
  NOR2_X1 U88 ( .A1(n305), .A2(n306), .ZN(n286) );
  AOI21_X1 U89 ( .B1(n289), .B2(n142), .A(n290), .ZN(n288) );
  NAND2_X1 U90 ( .A1(n146), .A2(n292), .ZN(n154) );
  NAND2_X1 U91 ( .A1(n82), .A2(n237), .ZN(n96) );
  NAND2_X1 U92 ( .A1(n30), .A2(n175), .ZN(n38) );
  NAND2_X1 U93 ( .A1(n119), .A2(n263), .ZN(n130) );
  NAND2_X1 U94 ( .A1(n39), .A2(n183), .ZN(n41) );
  NAND2_X1 U95 ( .A1(n97), .A2(n245), .ZN(n99) );
  INV_X1 U96 ( .A(n68), .ZN(n834) );
  NAND2_X1 U97 ( .A1(n131), .A2(n276), .ZN(n133) );
  INV_X1 U98 ( .A(n149), .ZN(n866) );
  NAND2_X1 U99 ( .A1(n89), .A2(n69), .ZN(n88) );
  INV_X1 U100 ( .A(n89), .ZN(n838) );
  INV_X1 U101 ( .A(n198), .ZN(n833) );
  INV_X1 U102 ( .A(n86), .ZN(n843) );
  NAND2_X1 U103 ( .A1(n61), .A2(n204), .ZN(n55) );
  NAND2_X1 U104 ( .A1(n69), .A2(n216), .ZN(n72) );
  NOR2_X1 U105 ( .A1(n200), .A2(n201), .ZN(n193) );
  NAND2_X1 U106 ( .A1(n183), .A2(n204), .ZN(n200) );
  NAND2_X1 U107 ( .A1(n46), .A2(n45), .ZN(n201) );
  NAND2_X1 U108 ( .A1(n39), .A2(n40), .ZN(n36) );
  INV_X1 U109 ( .A(n56), .ZN(n829) );
  NAND2_X1 U110 ( .A1(n97), .A2(n98), .ZN(n94) );
  INV_X1 U111 ( .A(n106), .ZN(n845) );
  NAND2_X1 U112 ( .A1(n132), .A2(n131), .ZN(n135) );
  NAND2_X1 U113 ( .A1(n131), .A2(n132), .ZN(n128) );
  AND2_X1 U114 ( .A1(n59), .A2(n198), .ZN(n1) );
  NAND2_X1 U115 ( .A1(n70), .A2(n66), .ZN(n228) );
  NAND2_X1 U116 ( .A1(n136), .A2(n134), .ZN(n306) );
  NAND2_X1 U117 ( .A1(n276), .A2(n298), .ZN(n305) );
  INV_X1 U118 ( .A(n82), .ZN(n846) );
  NAND2_X1 U119 ( .A1(n257), .A2(n258), .ZN(n256) );
  NAND2_X1 U120 ( .A1(n858), .A2(n855), .ZN(n258) );
  INV_X1 U121 ( .A(n118), .ZN(n858) );
  INV_X1 U122 ( .A(n90), .ZN(n840) );
  INV_X1 U123 ( .A(n27), .ZN(n815) );
  NAND2_X1 U124 ( .A1(n225), .A2(n226), .ZN(n207) );
  NOR2_X1 U125 ( .A1(n227), .A2(n228), .ZN(n226) );
  AOI21_X1 U126 ( .B1(n233), .B2(n841), .A(n234), .ZN(n225) );
  NAND2_X1 U127 ( .A1(n216), .A2(n231), .ZN(n227) );
  NAND2_X1 U128 ( .A1(n147), .A2(n148), .ZN(n122) );
  AND2_X1 U129 ( .A1(n150), .A2(n6), .ZN(n148) );
  AND2_X1 U130 ( .A1(n149), .A2(n131), .ZN(n6) );
  INV_X1 U131 ( .A(n105), .ZN(n849) );
  AND2_X1 U132 ( .A1(n313), .A2(n98), .ZN(n112) );
  OR2_X1 U133 ( .A1(n115), .A2(n116), .ZN(n313) );
  AND2_X1 U134 ( .A1(n5), .A2(n15), .ZN(n165) );
  AND2_X1 U135 ( .A1(n31), .A2(n17), .ZN(n5) );
  AND2_X1 U136 ( .A1(n40), .A2(n27), .ZN(n179) );
  AND2_X1 U137 ( .A1(n98), .A2(n86), .ZN(n241) );
  INV_X1 U138 ( .A(n29), .ZN(n817) );
  INV_X1 U139 ( .A(n30), .ZN(n818) );
  OR2_X1 U140 ( .A1(n58), .A2(n55), .ZN(n194) );
  INV_X1 U141 ( .A(n146), .ZN(n872) );
  INV_X1 U142 ( .A(n9), .ZN(GE) );
  INV_X1 U143 ( .A(n263), .ZN(n862) );
  INV_X1 U144 ( .A(n175), .ZN(n820) );
  XNOR2_X1 U145 ( .A(B[31]), .B(A[31]), .ZN(n15) );
  NAND2_X1 U146 ( .A1(A[18]), .A2(n837), .ZN(n69) );
  INV_X1 U147 ( .A(B[18]), .ZN(n837) );
  NAND2_X1 U148 ( .A1(A[24]), .A2(n823), .ZN(n39) );
  INV_X1 U149 ( .A(B[24]), .ZN(n823) );
  NAND2_X1 U150 ( .A1(A[25]), .A2(n821), .ZN(n40) );
  INV_X1 U151 ( .A(B[25]), .ZN(n821) );
  NAND2_X1 U152 ( .A1(A[12]), .A2(n851), .ZN(n97) );
  INV_X1 U153 ( .A(B[12]), .ZN(n851) );
  NAND2_X1 U154 ( .A1(A[13]), .A2(n848), .ZN(n98) );
  INV_X1 U155 ( .A(B[13]), .ZN(n848) );
  NAND2_X1 U156 ( .A1(A[19]), .A2(n835), .ZN(n68) );
  INV_X1 U157 ( .A(B[19]), .ZN(n835) );
  XNOR2_X1 U158 ( .A(B[30]), .B(A[30]), .ZN(n17) );
  NAND2_X1 U159 ( .A1(A[6]), .A2(n865), .ZN(n131) );
  INV_X1 U160 ( .A(B[6]), .ZN(n865) );
  NAND2_X1 U161 ( .A1(A[27]), .A2(n816), .ZN(n27) );
  INV_X1 U162 ( .A(B[27]), .ZN(n816) );
  NOR2_X1 U163 ( .A1(B[31]), .A2(n876), .ZN(n13) );
  NAND2_X1 U164 ( .A1(A[26]), .A2(n819), .ZN(n30) );
  INV_X1 U165 ( .A(B[26]), .ZN(n819) );
  NAND2_X1 U166 ( .A1(A[17]), .A2(n839), .ZN(n89) );
  INV_X1 U167 ( .A(B[17]), .ZN(n839) );
  NAND2_X1 U168 ( .A1(A[7]), .A2(n863), .ZN(n132) );
  INV_X1 U169 ( .A(B[7]), .ZN(n863) );
  NAND2_X1 U170 ( .A1(A[8]), .A2(n861), .ZN(n119) );
  INV_X1 U171 ( .A(B[8]), .ZN(n861) );
  NAND2_X1 U172 ( .A1(A[16]), .A2(n842), .ZN(n90) );
  INV_X1 U173 ( .A(B[16]), .ZN(n842) );
  NAND2_X1 U174 ( .A1(A[14]), .A2(n847), .ZN(n82) );
  INV_X1 U175 ( .A(B[14]), .ZN(n847) );
  NAND2_X1 U176 ( .A1(A[15]), .A2(n844), .ZN(n86) );
  INV_X1 U177 ( .A(B[15]), .ZN(n844) );
  NAND2_X1 U178 ( .A1(A[9]), .A2(n857), .ZN(n116) );
  INV_X1 U179 ( .A(B[9]), .ZN(n857) );
  NAND2_X1 U180 ( .A1(A[23]), .A2(n825), .ZN(n60) );
  INV_X1 U181 ( .A(B[23]), .ZN(n825) );
  NAND2_X1 U182 ( .A1(A[28]), .A2(n814), .ZN(n32) );
  INV_X1 U183 ( .A(B[28]), .ZN(n814) );
  NAND2_X1 U184 ( .A1(A[22]), .A2(n828), .ZN(n61) );
  INV_X1 U185 ( .A(B[22]), .ZN(n828) );
  NAND2_X1 U186 ( .A1(A[3]), .A2(n871), .ZN(n142) );
  INV_X1 U187 ( .A(B[3]), .ZN(n871) );
  NAND2_X1 U188 ( .A1(A[20]), .A2(n832), .ZN(n59) );
  INV_X1 U189 ( .A(B[20]), .ZN(n832) );
  NAND2_X1 U190 ( .A1(A[21]), .A2(n830), .ZN(n56) );
  INV_X1 U191 ( .A(B[21]), .ZN(n830) );
  NAND2_X1 U192 ( .A1(A[11]), .A2(n853), .ZN(n120) );
  INV_X1 U193 ( .A(B[11]), .ZN(n853) );
  NAND2_X1 U194 ( .A1(B[12]), .A2(n895), .ZN(n245) );
  INV_X1 U195 ( .A(A[12]), .ZN(n895) );
  NAND2_X1 U196 ( .A1(A[10]), .A2(n856), .ZN(n121) );
  INV_X1 U197 ( .A(B[10]), .ZN(n856) );
  NAND2_X1 U198 ( .A1(A[29]), .A2(n812), .ZN(n31) );
  INV_X1 U199 ( .A(B[29]), .ZN(n812) );
  NAND2_X1 U200 ( .A1(B[24]), .A2(n883), .ZN(n183) );
  INV_X1 U201 ( .A(A[24]), .ZN(n883) );
  NAND2_X1 U202 ( .A1(B[18]), .A2(n889), .ZN(n216) );
  INV_X1 U203 ( .A(A[18]), .ZN(n889) );
  NAND2_X1 U204 ( .A1(B[7]), .A2(n900), .ZN(n136) );
  INV_X1 U205 ( .A(A[7]), .ZN(n900) );
  NAND2_X1 U206 ( .A1(B[6]), .A2(n901), .ZN(n276) );
  INV_X1 U207 ( .A(A[6]), .ZN(n901) );
  NAND2_X1 U208 ( .A1(B[13]), .A2(n894), .ZN(n105) );
  INV_X1 U209 ( .A(A[13]), .ZN(n894) );
  NAND2_X1 U210 ( .A1(B[19]), .A2(n888), .ZN(n70) );
  INV_X1 U211 ( .A(A[19]), .ZN(n888) );
  NAND2_X1 U212 ( .A1(A[2]), .A2(n873), .ZN(n146) );
  INV_X1 U213 ( .A(B[2]), .ZN(n873) );
  NAND2_X1 U214 ( .A1(B[9]), .A2(n898), .ZN(n118) );
  INV_X1 U215 ( .A(A[9]), .ZN(n898) );
  NAND2_X1 U216 ( .A1(B[25]), .A2(n882), .ZN(n46) );
  INV_X1 U217 ( .A(A[25]), .ZN(n882) );
  NAND2_X1 U218 ( .A1(A[5]), .A2(n867), .ZN(n149) );
  INV_X1 U219 ( .A(B[5]), .ZN(n867) );
  NAND2_X1 U220 ( .A1(B[10]), .A2(n897), .ZN(n264) );
  INV_X1 U221 ( .A(A[10]), .ZN(n897) );
  NAND2_X1 U222 ( .A1(A[4]), .A2(n869), .ZN(n150) );
  INV_X1 U223 ( .A(B[4]), .ZN(n869) );
  NAND2_X1 U224 ( .A1(B[8]), .A2(n899), .ZN(n263) );
  INV_X1 U225 ( .A(A[8]), .ZN(n899) );
  INV_X1 U226 ( .A(A[31]), .ZN(n876) );
  NAND2_X1 U227 ( .A1(B[21]), .A2(n886), .ZN(n58) );
  INV_X1 U228 ( .A(A[21]), .ZN(n886) );
  NAND2_X1 U229 ( .A1(B[11]), .A2(n896), .ZN(n103) );
  INV_X1 U230 ( .A(A[11]), .ZN(n896) );
  NAND2_X1 U231 ( .A1(B[22]), .A2(n885), .ZN(n204) );
  INV_X1 U232 ( .A(A[22]), .ZN(n885) );
  INV_X1 U233 ( .A(A[1]), .ZN(n906) );
  NAND2_X1 U234 ( .A1(B[16]), .A2(n891), .ZN(n231) );
  INV_X1 U235 ( .A(A[16]), .ZN(n891) );
  NAND2_X1 U236 ( .A1(B[14]), .A2(n893), .ZN(n237) );
  INV_X1 U237 ( .A(A[14]), .ZN(n893) );
  NAND2_X1 U238 ( .A1(B[23]), .A2(n884), .ZN(n45) );
  INV_X1 U239 ( .A(A[23]), .ZN(n884) );
  NAND2_X1 U240 ( .A1(B[17]), .A2(n890), .ZN(n66) );
  INV_X1 U241 ( .A(A[17]), .ZN(n890) );
  NAND2_X1 U242 ( .A1(B[15]), .A2(n892), .ZN(n106) );
  INV_X1 U243 ( .A(A[15]), .ZN(n892) );
  NAND2_X1 U244 ( .A1(B[3]), .A2(n904), .ZN(n144) );
  INV_X1 U245 ( .A(A[3]), .ZN(n904) );
  NAND2_X1 U246 ( .A1(B[27]), .A2(n880), .ZN(n29) );
  INV_X1 U247 ( .A(A[27]), .ZN(n880) );
  NAND2_X1 U248 ( .A1(B[26]), .A2(n881), .ZN(n175) );
  INV_X1 U249 ( .A(A[26]), .ZN(n881) );
  NAND2_X1 U250 ( .A1(B[4]), .A2(n903), .ZN(n298) );
  INV_X1 U251 ( .A(A[4]), .ZN(n903) );
  NAND2_X1 U252 ( .A1(B[2]), .A2(n905), .ZN(n292) );
  INV_X1 U253 ( .A(A[2]), .ZN(n905) );
  NAND2_X1 U254 ( .A1(B[20]), .A2(n887), .ZN(n198) );
  INV_X1 U255 ( .A(A[20]), .ZN(n887) );
  INV_X1 U256 ( .A(A[30]), .ZN(n877) );
  NAND2_X1 U257 ( .A1(n161), .A2(n162), .ZN(n9) );
  NOR2_X1 U258 ( .A1(n4), .A2(n7), .ZN(n161) );
  OAI21_X1 U259 ( .B1(n163), .B2(n164), .A(n165), .ZN(n162) );
  AND3_X1 U260 ( .A1(B[30]), .A2(n877), .A3(n15), .ZN(n7) );
  NAND2_X1 U261 ( .A1(B[5]), .A2(n902), .ZN(n134) );
  INV_X1 U262 ( .A(A[5]), .ZN(n902) );
  NAND2_X1 U263 ( .A1(B[28]), .A2(n879), .ZN(n172) );
  INV_X1 U264 ( .A(A[28]), .ZN(n879) );
  NAND2_X1 U265 ( .A1(B[29]), .A2(n878), .ZN(n16) );
  INV_X1 U266 ( .A(A[29]), .ZN(n878) );
  INV_X1 U267 ( .A(B[1]), .ZN(n874) );
  AND3_X1 U268 ( .A1(A[30]), .A2(n811), .A3(n15), .ZN(n3) );
  INV_X1 U269 ( .A(B[30]), .ZN(n811) );
  AND2_X1 U270 ( .A1(B[31]), .A2(n876), .ZN(n4) );
  NAND2_X1 U271 ( .A1(n155), .A2(n156), .ZN(n152) );
  NAND2_X1 U272 ( .A1(A[0]), .A2(n875), .ZN(n156) );
  NAND2_X1 U273 ( .A1(A[1]), .A2(n874), .ZN(n155) );
  INV_X1 U274 ( .A(B[0]), .ZN(n875) );
  NAND2_X1 U275 ( .A1(n300), .A2(n301), .ZN(n294) );
  NAND2_X1 U276 ( .A1(B[1]), .A2(n906), .ZN(n300) );
  NAND2_X1 U277 ( .A1(B[0]), .A2(n907), .ZN(n301) );
  INV_X1 U278 ( .A(A[0]), .ZN(n907) );
  AND2_X1 U279 ( .A1(n303), .A2(n142), .ZN(n293) );
  NAND2_X1 U280 ( .A1(A[1]), .A2(n874), .ZN(n303) );
  AND2_X1 U290 ( .A1(n159), .A2(n144), .ZN(n151) );
  NAND2_X1 U291 ( .A1(B[1]), .A2(n906), .ZN(n159) );
endmodule


module COMPARATOR_M32 ( A, B, sel, OUTPUT );
  input [31:0] A;
  input [31:0] B;
  input [1:0] sel;
  output [31:0] OUTPUT;
  wire   N12, N15, N16, n5, n6, n16, n17;
  assign OUTPUT[1] = 1'b0;
  assign OUTPUT[2] = 1'b0;
  assign OUTPUT[3] = 1'b0;
  assign OUTPUT[4] = 1'b0;
  assign OUTPUT[5] = 1'b0;
  assign OUTPUT[6] = 1'b0;
  assign OUTPUT[7] = 1'b0;
  assign OUTPUT[8] = 1'b0;
  assign OUTPUT[9] = 1'b0;
  assign OUTPUT[10] = 1'b0;
  assign OUTPUT[11] = 1'b0;
  assign OUTPUT[12] = 1'b0;
  assign OUTPUT[13] = 1'b0;
  assign OUTPUT[14] = 1'b0;
  assign OUTPUT[15] = 1'b0;
  assign OUTPUT[16] = 1'b0;
  assign OUTPUT[17] = 1'b0;
  assign OUTPUT[18] = 1'b0;
  assign OUTPUT[19] = 1'b0;
  assign OUTPUT[20] = 1'b0;
  assign OUTPUT[21] = 1'b0;
  assign OUTPUT[22] = 1'b0;
  assign OUTPUT[23] = 1'b0;
  assign OUTPUT[24] = 1'b0;
  assign OUTPUT[25] = 1'b0;
  assign OUTPUT[26] = 1'b0;
  assign OUTPUT[27] = 1'b0;
  assign OUTPUT[28] = 1'b0;
  assign OUTPUT[29] = 1'b0;
  assign OUTPUT[30] = 1'b0;
  assign OUTPUT[31] = 1'b0;

  XOR2_X1 U8 ( .A(n16), .B(N12), .Z(n6) );
  COMPARATOR_M32_DW01_cmp6_1 r61 ( .A(A), .B(B), .TC(1'b0), .EQ(N12), .LE(N16), 
        .GE(N15) );
  INV_X1 U2 ( .A(sel[0]), .ZN(n16) );
  OAI22_X1 U4 ( .A1(n5), .A2(n17), .B1(sel[1]), .B2(n6), .ZN(OUTPUT[0]) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n17) );
  AOI22_X1 U6 ( .A1(N15), .A2(n16), .B1(N16), .B2(sel[0]), .ZN(n5) );
endmodule


module ALU_M32_C4 ( CODE, DATA1, DATA2, OUTALU );
  input [3:0] CODE;
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTALU;
  wire   \Comparison[1] , \COMPARATORout[0] , n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405;
  wire   [31:0] SHIFTERout;
  wire   [31:0] ADDERout;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  XOR2_X1 U209 ( .A(CODE[1]), .B(CODE[0]), .Z(n176) );
  SHIFTER_M32_N5 SHIFTOP ( .A(DATA1), .B(DATA2), .LEFT_RIGHT(CODE[0]), 
        .OUTPUT(SHIFTERout) );
  P4ADDER_n_bit32 ADDSUBOP ( .A(DATA1), .B(DATA2), .cin0(n1337), .S(ADDERout)
         );
  COMPARATOR_M32 COMPOP ( .A(DATA1), .B(DATA2), .sel({\Comparison[1] , n1405}), 
        .OUTPUT({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, \COMPARATORout[0] }) );
  NOR3_X1 U2 ( .A1(n1405), .A2(CODE[0]), .A3(n174), .ZN(n77) );
  BUF_X1 U3 ( .A(n75), .Z(n1326) );
  BUF_X1 U4 ( .A(n75), .Z(n1327) );
  BUF_X1 U5 ( .A(n75), .Z(n1328) );
  BUF_X1 U6 ( .A(n75), .Z(n1329) );
  BUF_X1 U7 ( .A(n77), .Z(n1317) );
  BUF_X1 U8 ( .A(n77), .Z(n1316) );
  BUF_X1 U9 ( .A(n77), .Z(n1319) );
  BUF_X1 U10 ( .A(n77), .Z(n1320) );
  BUF_X1 U11 ( .A(n77), .Z(n1318) );
  BUF_X1 U12 ( .A(n75), .Z(n1325) );
  AOI21_X1 U13 ( .B1(n1330), .B2(n1370), .A(n1321), .ZN(n170) );
  AOI221_X1 U14 ( .B1(n1327), .B2(n1402), .C1(DATA1[0]), .C2(n1322), .A(n1318), 
        .ZN(n171) );
  NOR2_X1 U15 ( .A1(n174), .A2(n173), .ZN(n75) );
  BUF_X1 U16 ( .A(n76), .Z(n1322) );
  BUF_X1 U17 ( .A(n76), .Z(n1323) );
  BUF_X1 U18 ( .A(n73), .Z(n1335) );
  BUF_X1 U19 ( .A(n73), .Z(n1334) );
  BUF_X1 U20 ( .A(n74), .Z(n1331) );
  BUF_X1 U21 ( .A(n74), .Z(n1332) );
  OAI221_X1 U22 ( .B1(n99), .B2(n1372), .C1(n100), .C2(n1340), .A(n101), .ZN(
        OUTALU[30]) );
  AOI21_X1 U23 ( .B1(n1329), .B2(n1340), .A(n1320), .ZN(n99) );
  AOI22_X1 U24 ( .A1(SHIFTERout[30]), .A2(n1334), .B1(ADDERout[30]), .B2(n1332), .ZN(n101) );
  AOI221_X1 U25 ( .B1(n1325), .B2(n1372), .C1(DATA1[30]), .C2(n1323), .A(n1316), .ZN(n100) );
  OAI221_X1 U26 ( .B1(n78), .B2(n1394), .C1(n79), .C2(n1362), .A(n80), .ZN(
        OUTALU[8]) );
  AOI21_X1 U27 ( .B1(n1330), .B2(n1362), .A(n1320), .ZN(n78) );
  AOI22_X1 U28 ( .A1(SHIFTERout[8]), .A2(n1334), .B1(ADDERout[8]), .B2(n1333), 
        .ZN(n80) );
  AOI221_X1 U29 ( .B1(n1325), .B2(n1394), .C1(DATA1[8]), .C2(n1324), .A(n1316), 
        .ZN(n79) );
  OAI221_X1 U30 ( .B1(n70), .B2(n1393), .C1(n71), .C2(n1361), .A(n72), .ZN(
        OUTALU[9]) );
  AOI21_X1 U31 ( .B1(n1330), .B2(n1361), .A(n1321), .ZN(n70) );
  AOI22_X1 U32 ( .A1(SHIFTERout[9]), .A2(n1334), .B1(ADDERout[9]), .B2(n1333), 
        .ZN(n72) );
  AOI221_X1 U33 ( .B1(n1326), .B2(n1393), .C1(n1324), .C2(DATA1[9]), .A(n1317), 
        .ZN(n71) );
  OAI221_X1 U34 ( .B1(n165), .B2(n1392), .C1(n166), .C2(n1360), .A(n167), .ZN(
        OUTALU[10]) );
  AOI21_X1 U35 ( .B1(n1330), .B2(n1360), .A(n1320), .ZN(n165) );
  AOI22_X1 U36 ( .A1(SHIFTERout[10]), .A2(n1336), .B1(ADDERout[10]), .B2(n1331), .ZN(n167) );
  AOI221_X1 U37 ( .B1(n1327), .B2(n1392), .C1(DATA1[10]), .C2(n1322), .A(n1318), .ZN(n166) );
  OAI221_X1 U38 ( .B1(n162), .B2(n1391), .C1(n163), .C2(n1359), .A(n164), .ZN(
        OUTALU[11]) );
  AOI21_X1 U39 ( .B1(n1329), .B2(n1359), .A(n1320), .ZN(n162) );
  AOI22_X1 U40 ( .A1(SHIFTERout[11]), .A2(n1336), .B1(ADDERout[11]), .B2(n1331), .ZN(n164) );
  AOI221_X1 U41 ( .B1(n1327), .B2(n1391), .C1(DATA1[11]), .C2(n1322), .A(n1318), .ZN(n163) );
  OAI221_X1 U42 ( .B1(n159), .B2(n1390), .C1(n160), .C2(n1358), .A(n161), .ZN(
        OUTALU[12]) );
  AOI21_X1 U43 ( .B1(n1329), .B2(n1358), .A(n1320), .ZN(n159) );
  AOI22_X1 U44 ( .A1(SHIFTERout[12]), .A2(n1336), .B1(ADDERout[12]), .B2(n1331), .ZN(n161) );
  AOI221_X1 U45 ( .B1(n1327), .B2(n1390), .C1(DATA1[12]), .C2(n1322), .A(n1318), .ZN(n160) );
  OAI221_X1 U46 ( .B1(n156), .B2(n1389), .C1(n157), .C2(n1357), .A(n158), .ZN(
        OUTALU[13]) );
  AOI21_X1 U47 ( .B1(n1329), .B2(n1357), .A(n1320), .ZN(n156) );
  AOI22_X1 U48 ( .A1(SHIFTERout[13]), .A2(n1336), .B1(ADDERout[13]), .B2(n1331), .ZN(n158) );
  AOI221_X1 U49 ( .B1(n1327), .B2(n1389), .C1(DATA1[13]), .C2(n1322), .A(n1318), .ZN(n157) );
  OAI221_X1 U50 ( .B1(n153), .B2(n1388), .C1(n154), .C2(n1356), .A(n155), .ZN(
        OUTALU[14]) );
  AOI21_X1 U51 ( .B1(n1328), .B2(n1356), .A(n1319), .ZN(n153) );
  AOI22_X1 U52 ( .A1(SHIFTERout[14]), .A2(n1336), .B1(ADDERout[14]), .B2(n1331), .ZN(n155) );
  AOI221_X1 U53 ( .B1(n1327), .B2(n1388), .C1(DATA1[14]), .C2(n1322), .A(n1318), .ZN(n154) );
  OAI221_X1 U54 ( .B1(n150), .B2(n1387), .C1(n151), .C2(n1355), .A(n152), .ZN(
        OUTALU[15]) );
  AOI21_X1 U55 ( .B1(n1329), .B2(n1355), .A(n1319), .ZN(n150) );
  AOI22_X1 U56 ( .A1(SHIFTERout[15]), .A2(n1336), .B1(ADDERout[15]), .B2(n1331), .ZN(n152) );
  AOI221_X1 U57 ( .B1(n1327), .B2(n1387), .C1(DATA1[15]), .C2(n1322), .A(n1318), .ZN(n151) );
  OAI221_X1 U58 ( .B1(n147), .B2(n1386), .C1(n148), .C2(n1354), .A(n149), .ZN(
        OUTALU[16]) );
  AOI21_X1 U59 ( .B1(n1328), .B2(n1354), .A(n1319), .ZN(n147) );
  AOI22_X1 U60 ( .A1(SHIFTERout[16]), .A2(n1336), .B1(ADDERout[16]), .B2(n1331), .ZN(n149) );
  AOI221_X1 U61 ( .B1(n1326), .B2(n1386), .C1(DATA1[16]), .C2(n1322), .A(n1317), .ZN(n148) );
  OAI221_X1 U62 ( .B1(n144), .B2(n1385), .C1(n145), .C2(n1353), .A(n146), .ZN(
        OUTALU[17]) );
  AOI21_X1 U63 ( .B1(n1328), .B2(n1353), .A(n1319), .ZN(n144) );
  AOI22_X1 U64 ( .A1(SHIFTERout[17]), .A2(n1335), .B1(ADDERout[17]), .B2(n1331), .ZN(n146) );
  AOI221_X1 U65 ( .B1(n1327), .B2(n1385), .C1(DATA1[17]), .C2(n1322), .A(n1318), .ZN(n145) );
  OAI221_X1 U66 ( .B1(n141), .B2(n1384), .C1(n142), .C2(n1352), .A(n143), .ZN(
        OUTALU[18]) );
  AOI21_X1 U67 ( .B1(n1328), .B2(n1352), .A(n1319), .ZN(n141) );
  AOI22_X1 U68 ( .A1(SHIFTERout[18]), .A2(n1335), .B1(ADDERout[18]), .B2(n1331), .ZN(n143) );
  AOI221_X1 U69 ( .B1(n1326), .B2(n1384), .C1(DATA1[18]), .C2(n1322), .A(n1317), .ZN(n142) );
  OAI221_X1 U70 ( .B1(n138), .B2(n1383), .C1(n139), .C2(n1351), .A(n140), .ZN(
        OUTALU[19]) );
  AOI21_X1 U71 ( .B1(n1327), .B2(n1351), .A(n1318), .ZN(n138) );
  AOI22_X1 U72 ( .A1(SHIFTERout[19]), .A2(n1335), .B1(ADDERout[19]), .B2(n1331), .ZN(n140) );
  AOI221_X1 U73 ( .B1(n1326), .B2(n1383), .C1(DATA1[19]), .C2(n1322), .A(n1317), .ZN(n139) );
  OAI221_X1 U74 ( .B1(n132), .B2(n1382), .C1(n133), .C2(n1350), .A(n134), .ZN(
        OUTALU[20]) );
  AOI21_X1 U75 ( .B1(n1328), .B2(n1350), .A(n1319), .ZN(n132) );
  AOI22_X1 U76 ( .A1(SHIFTERout[20]), .A2(n1335), .B1(ADDERout[20]), .B2(n1332), .ZN(n134) );
  AOI221_X1 U77 ( .B1(n1326), .B2(n1382), .C1(DATA1[20]), .C2(n1323), .A(n1317), .ZN(n133) );
  OAI221_X1 U78 ( .B1(n129), .B2(n1381), .C1(n130), .C2(n1349), .A(n131), .ZN(
        OUTALU[21]) );
  AOI21_X1 U79 ( .B1(n1327), .B2(n1349), .A(n1318), .ZN(n129) );
  AOI22_X1 U80 ( .A1(SHIFTERout[21]), .A2(n1335), .B1(ADDERout[21]), .B2(n1332), .ZN(n131) );
  AOI221_X1 U81 ( .B1(n1326), .B2(n1381), .C1(DATA1[21]), .C2(n1323), .A(n1317), .ZN(n130) );
  OAI221_X1 U82 ( .B1(n126), .B2(n1380), .C1(n127), .C2(n1348), .A(n128), .ZN(
        OUTALU[22]) );
  AOI21_X1 U83 ( .B1(n1327), .B2(n1348), .A(n1318), .ZN(n126) );
  AOI22_X1 U84 ( .A1(SHIFTERout[22]), .A2(n1335), .B1(ADDERout[22]), .B2(n1332), .ZN(n128) );
  AOI221_X1 U85 ( .B1(n1326), .B2(n1380), .C1(DATA1[22]), .C2(n1323), .A(n1317), .ZN(n127) );
  OAI221_X1 U86 ( .B1(n123), .B2(n1379), .C1(n124), .C2(n1347), .A(n125), .ZN(
        OUTALU[23]) );
  AOI21_X1 U87 ( .B1(n1328), .B2(n1347), .A(n1319), .ZN(n123) );
  AOI22_X1 U88 ( .A1(SHIFTERout[23]), .A2(n1335), .B1(ADDERout[23]), .B2(n1332), .ZN(n125) );
  AOI221_X1 U89 ( .B1(n1326), .B2(n1379), .C1(DATA1[23]), .C2(n1323), .A(n1317), .ZN(n124) );
  OAI221_X1 U90 ( .B1(n120), .B2(n1378), .C1(n121), .C2(n1346), .A(n122), .ZN(
        OUTALU[24]) );
  AOI21_X1 U91 ( .B1(n1328), .B2(n1346), .A(n1319), .ZN(n120) );
  AOI22_X1 U92 ( .A1(SHIFTERout[24]), .A2(n1335), .B1(ADDERout[24]), .B2(n1332), .ZN(n122) );
  AOI221_X1 U93 ( .B1(n1326), .B2(n1378), .C1(DATA1[24]), .C2(n1323), .A(n1317), .ZN(n121) );
  OAI221_X1 U94 ( .B1(n117), .B2(n1377), .C1(n118), .C2(n1345), .A(n119), .ZN(
        OUTALU[25]) );
  AOI21_X1 U95 ( .B1(n1328), .B2(n1345), .A(n1319), .ZN(n117) );
  AOI22_X1 U96 ( .A1(SHIFTERout[25]), .A2(n1335), .B1(ADDERout[25]), .B2(n1332), .ZN(n119) );
  AOI221_X1 U97 ( .B1(n1326), .B2(n1377), .C1(DATA1[25]), .C2(n1323), .A(n1317), .ZN(n118) );
  OAI221_X1 U98 ( .B1(n114), .B2(n1376), .C1(n115), .C2(n1344), .A(n116), .ZN(
        OUTALU[26]) );
  AOI21_X1 U99 ( .B1(n1328), .B2(n1344), .A(n1319), .ZN(n114) );
  AOI22_X1 U100 ( .A1(SHIFTERout[26]), .A2(n1335), .B1(ADDERout[26]), .B2(
        n1332), .ZN(n116) );
  AOI221_X1 U101 ( .B1(n1326), .B2(n1376), .C1(DATA1[26]), .C2(n1323), .A(
        n1317), .ZN(n115) );
  OAI221_X1 U102 ( .B1(n111), .B2(n1375), .C1(n112), .C2(n1343), .A(n113), 
        .ZN(OUTALU[27]) );
  AOI21_X1 U103 ( .B1(n1328), .B2(n1343), .A(n1319), .ZN(n111) );
  AOI22_X1 U104 ( .A1(SHIFTERout[27]), .A2(n1335), .B1(ADDERout[27]), .B2(
        n1332), .ZN(n113) );
  AOI221_X1 U105 ( .B1(n1325), .B2(n1375), .C1(DATA1[27]), .C2(n1323), .A(
        n1316), .ZN(n112) );
  OAI221_X1 U106 ( .B1(n108), .B2(n1374), .C1(n109), .C2(n1342), .A(n110), 
        .ZN(OUTALU[28]) );
  AOI21_X1 U107 ( .B1(n1328), .B2(n1342), .A(n1319), .ZN(n108) );
  AOI22_X1 U108 ( .A1(SHIFTERout[28]), .A2(n1334), .B1(ADDERout[28]), .B2(
        n1332), .ZN(n110) );
  AOI221_X1 U109 ( .B1(n1325), .B2(n1374), .C1(DATA1[28]), .C2(n1323), .A(
        n1316), .ZN(n109) );
  OAI221_X1 U110 ( .B1(n105), .B2(n1373), .C1(n106), .C2(n1341), .A(n107), 
        .ZN(OUTALU[29]) );
  AOI21_X1 U111 ( .B1(n1329), .B2(n1341), .A(n1320), .ZN(n105) );
  AOI22_X1 U112 ( .A1(SHIFTERout[29]), .A2(n1334), .B1(ADDERout[29]), .B2(
        n1332), .ZN(n107) );
  AOI221_X1 U113 ( .B1(n1325), .B2(n1373), .C1(DATA1[29]), .C2(n1323), .A(
        n1316), .ZN(n106) );
  OAI221_X1 U114 ( .B1(n96), .B2(n1371), .C1(n97), .C2(n1339), .A(n98), .ZN(
        OUTALU[31]) );
  AOI21_X1 U115 ( .B1(n1329), .B2(n1339), .A(n1320), .ZN(n96) );
  AOI22_X1 U116 ( .A1(SHIFTERout[31]), .A2(n1334), .B1(ADDERout[31]), .B2(
        n1333), .ZN(n98) );
  AOI221_X1 U117 ( .B1(n1325), .B2(n1371), .C1(DATA1[31]), .C2(n1324), .A(
        n1316), .ZN(n97) );
  BUF_X1 U118 ( .A(n76), .Z(n1324) );
  BUF_X1 U119 ( .A(n74), .Z(n1333) );
  BUF_X1 U120 ( .A(n73), .Z(n1336) );
  INV_X1 U121 ( .A(DATA2[31]), .ZN(n1339) );
  INV_X1 U122 ( .A(DATA1[30]), .ZN(n1372) );
  NAND2_X1 U123 ( .A1(n1405), .A2(n1337), .ZN(\Comparison[1] ) );
  INV_X1 U124 ( .A(DATA1[29]), .ZN(n1373) );
  INV_X1 U125 ( .A(DATA1[25]), .ZN(n1377) );
  INV_X1 U126 ( .A(DATA1[15]), .ZN(n1387) );
  INV_X1 U127 ( .A(DATA1[24]), .ZN(n1378) );
  INV_X1 U128 ( .A(DATA1[31]), .ZN(n1371) );
  INV_X1 U129 ( .A(DATA1[13]), .ZN(n1389) );
  INV_X1 U130 ( .A(DATA1[22]), .ZN(n1380) );
  INV_X1 U131 ( .A(DATA1[28]), .ZN(n1374) );
  INV_X1 U132 ( .A(DATA1[12]), .ZN(n1390) );
  INV_X1 U133 ( .A(DATA1[23]), .ZN(n1379) );
  INV_X1 U134 ( .A(DATA1[26]), .ZN(n1376) );
  INV_X1 U135 ( .A(DATA1[17]), .ZN(n1385) );
  INV_X1 U136 ( .A(DATA1[9]), .ZN(n1393) );
  INV_X1 U137 ( .A(DATA1[8]), .ZN(n1394) );
  INV_X1 U138 ( .A(DATA1[16]), .ZN(n1386) );
  INV_X1 U139 ( .A(DATA1[20]), .ZN(n1382) );
  INV_X1 U140 ( .A(DATA1[11]), .ZN(n1391) );
  INV_X1 U141 ( .A(DATA1[19]), .ZN(n1383) );
  INV_X1 U142 ( .A(DATA1[27]), .ZN(n1375) );
  INV_X1 U143 ( .A(DATA1[10]), .ZN(n1392) );
  INV_X1 U144 ( .A(DATA1[14]), .ZN(n1388) );
  INV_X1 U145 ( .A(DATA1[18]), .ZN(n1384) );
  INV_X1 U146 ( .A(DATA1[21]), .ZN(n1381) );
  INV_X1 U147 ( .A(DATA1[1]), .ZN(n1401) );
  INV_X1 U148 ( .A(DATA1[2]), .ZN(n1400) );
  INV_X1 U149 ( .A(DATA1[4]), .ZN(n1398) );
  INV_X1 U150 ( .A(DATA1[5]), .ZN(n1397) );
  INV_X1 U151 ( .A(DATA1[6]), .ZN(n1396) );
  INV_X1 U152 ( .A(DATA1[3]), .ZN(n1399) );
  INV_X1 U153 ( .A(DATA1[7]), .ZN(n1395) );
  INV_X1 U154 ( .A(DATA1[0]), .ZN(n1402) );
  INV_X1 U155 ( .A(DATA2[9]), .ZN(n1361) );
  INV_X1 U156 ( .A(DATA2[8]), .ZN(n1362) );
  INV_X1 U157 ( .A(DATA2[13]), .ZN(n1357) );
  INV_X1 U158 ( .A(DATA2[7]), .ZN(n1363) );
  INV_X1 U159 ( .A(DATA2[10]), .ZN(n1360) );
  INV_X1 U160 ( .A(DATA2[12]), .ZN(n1358) );
  INV_X1 U161 ( .A(DATA2[11]), .ZN(n1359) );
  INV_X1 U162 ( .A(DATA2[30]), .ZN(n1340) );
  INV_X1 U163 ( .A(DATA2[21]), .ZN(n1349) );
  INV_X1 U164 ( .A(DATA2[20]), .ZN(n1350) );
  INV_X1 U165 ( .A(DATA2[22]), .ZN(n1348) );
  INV_X1 U166 ( .A(DATA2[29]), .ZN(n1341) );
  INV_X1 U167 ( .A(DATA2[17]), .ZN(n1353) );
  INV_X1 U168 ( .A(DATA2[23]), .ZN(n1347) );
  INV_X1 U169 ( .A(DATA2[19]), .ZN(n1351) );
  INV_X1 U170 ( .A(DATA2[18]), .ZN(n1352) );
  INV_X1 U171 ( .A(DATA2[16]), .ZN(n1354) );
  INV_X1 U172 ( .A(DATA2[28]), .ZN(n1342) );
  INV_X1 U173 ( .A(DATA2[15]), .ZN(n1355) );
  INV_X1 U174 ( .A(DATA2[14]), .ZN(n1356) );
  INV_X1 U175 ( .A(DATA2[25]), .ZN(n1345) );
  INV_X1 U176 ( .A(DATA2[24]), .ZN(n1346) );
  INV_X1 U177 ( .A(DATA2[0]), .ZN(n1370) );
  INV_X1 U178 ( .A(DATA2[27]), .ZN(n1343) );
  INV_X1 U179 ( .A(DATA2[26]), .ZN(n1344) );
  INV_X1 U180 ( .A(DATA2[6]), .ZN(n1364) );
  INV_X1 U181 ( .A(DATA2[1]), .ZN(n1369) );
  INV_X1 U182 ( .A(DATA2[5]), .ZN(n1365) );
  INV_X1 U183 ( .A(DATA2[2]), .ZN(n1368) );
  INV_X1 U184 ( .A(DATA2[3]), .ZN(n1367) );
  INV_X1 U185 ( .A(DATA2[4]), .ZN(n1366) );
  NOR3_X1 U186 ( .A1(n1337), .A2(CODE[1]), .A3(n174), .ZN(n76) );
  OAI21_X1 U187 ( .B1(\Comparison[1] ), .B2(n174), .A(n175), .ZN(n74) );
  OR3_X1 U188 ( .A1(CODE[2]), .A2(CODE[3]), .A3(n173), .ZN(n175) );
  OAI221_X1 U189 ( .B1(n135), .B2(n1401), .C1(n136), .C2(n1369), .A(n137), 
        .ZN(OUTALU[1]) );
  AOI21_X1 U190 ( .B1(n1327), .B2(n1369), .A(n1318), .ZN(n135) );
  AOI22_X1 U191 ( .A1(SHIFTERout[1]), .A2(n1335), .B1(ADDERout[1]), .B2(n1331), 
        .ZN(n137) );
  AOI221_X1 U192 ( .B1(n1326), .B2(n1401), .C1(DATA1[1]), .C2(n1322), .A(n1317), .ZN(n136) );
  OAI221_X1 U193 ( .B1(n102), .B2(n1400), .C1(n103), .C2(n1368), .A(n104), 
        .ZN(OUTALU[2]) );
  AOI21_X1 U194 ( .B1(n1328), .B2(n1368), .A(n1319), .ZN(n102) );
  AOI22_X1 U195 ( .A1(SHIFTERout[2]), .A2(n1334), .B1(ADDERout[2]), .B2(n1332), 
        .ZN(n104) );
  AOI221_X1 U196 ( .B1(n1325), .B2(n1400), .C1(DATA1[2]), .C2(n1323), .A(n1316), .ZN(n103) );
  OAI221_X1 U197 ( .B1(n93), .B2(n1399), .C1(n94), .C2(n1367), .A(n95), .ZN(
        OUTALU[3]) );
  AOI21_X1 U198 ( .B1(n1329), .B2(n1367), .A(n1320), .ZN(n93) );
  AOI22_X1 U199 ( .A1(SHIFTERout[3]), .A2(n1334), .B1(ADDERout[3]), .B2(n1333), 
        .ZN(n95) );
  AOI221_X1 U200 ( .B1(n1325), .B2(n1399), .C1(DATA1[3]), .C2(n1324), .A(n1316), .ZN(n94) );
  OAI221_X1 U201 ( .B1(n90), .B2(n1398), .C1(n91), .C2(n1366), .A(n92), .ZN(
        OUTALU[4]) );
  AOI21_X1 U202 ( .B1(n1329), .B2(n1366), .A(n1320), .ZN(n90) );
  AOI22_X1 U203 ( .A1(SHIFTERout[4]), .A2(n1334), .B1(ADDERout[4]), .B2(n1333), 
        .ZN(n92) );
  AOI221_X1 U204 ( .B1(n1325), .B2(n1398), .C1(DATA1[4]), .C2(n1324), .A(n1316), .ZN(n91) );
  OAI221_X1 U205 ( .B1(n87), .B2(n1397), .C1(n88), .C2(n1365), .A(n89), .ZN(
        OUTALU[5]) );
  AOI21_X1 U206 ( .B1(n1329), .B2(n1365), .A(n1320), .ZN(n87) );
  AOI22_X1 U207 ( .A1(SHIFTERout[5]), .A2(n1334), .B1(ADDERout[5]), .B2(n1333), 
        .ZN(n89) );
  AOI221_X1 U208 ( .B1(n1325), .B2(n1397), .C1(DATA1[5]), .C2(n1324), .A(n1316), .ZN(n88) );
  OAI221_X1 U210 ( .B1(n84), .B2(n1396), .C1(n85), .C2(n1364), .A(n86), .ZN(
        OUTALU[6]) );
  AOI21_X1 U211 ( .B1(n1329), .B2(n1364), .A(n1320), .ZN(n84) );
  AOI22_X1 U212 ( .A1(SHIFTERout[6]), .A2(n1334), .B1(ADDERout[6]), .B2(n1333), 
        .ZN(n86) );
  AOI221_X1 U213 ( .B1(n1325), .B2(n1396), .C1(DATA1[6]), .C2(n1324), .A(n1316), .ZN(n85) );
  OAI221_X1 U214 ( .B1(n81), .B2(n1395), .C1(n82), .C2(n1363), .A(n83), .ZN(
        OUTALU[7]) );
  AOI21_X1 U215 ( .B1(n1329), .B2(n1363), .A(n1320), .ZN(n81) );
  AOI22_X1 U216 ( .A1(SHIFTERout[7]), .A2(n1334), .B1(ADDERout[7]), .B2(n1333), 
        .ZN(n83) );
  AOI221_X1 U217 ( .B1(n1325), .B2(n1395), .C1(DATA1[7]), .C2(n1324), .A(n1316), .ZN(n82) );
  NAND2_X1 U218 ( .A1(CODE[2]), .A2(n1403), .ZN(n174) );
  INV_X1 U219 ( .A(CODE[1]), .ZN(n1405) );
  NAND4_X1 U220 ( .A1(\COMPARATORout[0] ), .A2(CODE[3]), .A3(n173), .A4(n1404), 
        .ZN(n172) );
  NAND2_X1 U221 ( .A1(CODE[0]), .A2(CODE[1]), .ZN(n173) );
  AND3_X1 U222 ( .A1(n1404), .A2(n1403), .A3(n176), .ZN(n73) );
  INV_X1 U223 ( .A(CODE[2]), .ZN(n1404) );
  INV_X1 U224 ( .A(CODE[3]), .ZN(n1403) );
  INV_X1 U225 ( .A(n168), .ZN(OUTALU[0]) );
  AOI221_X1 U226 ( .B1(SHIFTERout[0]), .B2(n1336), .C1(ADDERout[0]), .C2(n1331), .A(n169), .ZN(n168) );
  OAI221_X1 U227 ( .B1(n170), .B2(n1402), .C1(n171), .C2(n1370), .A(n172), 
        .ZN(n169) );
  CLKBUF_X1 U228 ( .A(n77), .Z(n1321) );
  CLKBUF_X1 U229 ( .A(n75), .Z(n1330) );
  INV_X1 U230 ( .A(CODE[0]), .ZN(n1337) );
endmodule


module reg_5 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n367), .Z(n329) );
  BUF_X1 U4 ( .A(n367), .Z(n328) );
  BUF_X1 U5 ( .A(n367), .Z(n330) );
  BUF_X1 U6 ( .A(n368), .Z(n331) );
  BUF_X1 U7 ( .A(n368), .Z(n332) );
  BUF_X1 U8 ( .A(n368), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n367) );
  OAI22_X1 U10 ( .A1(n333), .A2(n36), .B1(n330), .B2(n366), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n366) );
  OAI22_X1 U12 ( .A1(n333), .A2(n37), .B1(n330), .B2(n365), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n365) );
  OAI22_X1 U14 ( .A1(n333), .A2(n38), .B1(n330), .B2(n364), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n364) );
  OAI22_X1 U16 ( .A1(n333), .A2(n39), .B1(n330), .B2(n363), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n363) );
  OAI22_X1 U18 ( .A1(n333), .A2(n40), .B1(n330), .B2(n362), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n362) );
  OAI22_X1 U20 ( .A1(n333), .A2(n41), .B1(n330), .B2(n361), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n361) );
  OAI22_X1 U22 ( .A1(n333), .A2(n42), .B1(n330), .B2(n360), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n360) );
  OAI22_X1 U24 ( .A1(n332), .A2(n43), .B1(n330), .B2(n359), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n359) );
  OAI22_X1 U26 ( .A1(n332), .A2(n44), .B1(n329), .B2(n358), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n358) );
  OAI22_X1 U28 ( .A1(n332), .A2(n45), .B1(n329), .B2(n357), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n357) );
  OAI22_X1 U30 ( .A1(n332), .A2(n46), .B1(n329), .B2(n356), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n356) );
  OAI22_X1 U32 ( .A1(n332), .A2(n47), .B1(n329), .B2(n355), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n355) );
  OAI22_X1 U34 ( .A1(n332), .A2(n48), .B1(n329), .B2(n354), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n354) );
  OAI22_X1 U36 ( .A1(n332), .A2(n49), .B1(n329), .B2(n353), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n353) );
  OAI22_X1 U38 ( .A1(n332), .A2(n50), .B1(n329), .B2(n352), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n352) );
  OAI22_X1 U40 ( .A1(n332), .A2(n51), .B1(n329), .B2(n351), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n351) );
  OAI22_X1 U42 ( .A1(n332), .A2(n52), .B1(n329), .B2(n350), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n350) );
  OAI22_X1 U44 ( .A1(n332), .A2(n53), .B1(n329), .B2(n349), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n349) );
  OAI22_X1 U46 ( .A1(n332), .A2(n54), .B1(n329), .B2(n348), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n348) );
  OAI22_X1 U48 ( .A1(n332), .A2(n55), .B1(n329), .B2(n347), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n347) );
  OAI22_X1 U50 ( .A1(n331), .A2(n56), .B1(n328), .B2(n346), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n346) );
  OAI22_X1 U52 ( .A1(n331), .A2(n57), .B1(n328), .B2(n345), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n345) );
  OAI22_X1 U54 ( .A1(n331), .A2(n58), .B1(n328), .B2(n344), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n344) );
  OAI22_X1 U56 ( .A1(n331), .A2(n59), .B1(n328), .B2(n343), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n343) );
  OAI22_X1 U58 ( .A1(n331), .A2(n60), .B1(n328), .B2(n342), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n342) );
  OAI22_X1 U60 ( .A1(n331), .A2(n61), .B1(n328), .B2(n341), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n341) );
  OAI22_X1 U62 ( .A1(n331), .A2(n62), .B1(n328), .B2(n340), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n340) );
  OAI22_X1 U64 ( .A1(n331), .A2(n63), .B1(n328), .B2(n339), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n339) );
  OAI22_X1 U66 ( .A1(n331), .A2(n64), .B1(n328), .B2(n338), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n338) );
  OAI22_X1 U68 ( .A1(n331), .A2(n65), .B1(n328), .B2(n337), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n337) );
  OAI22_X1 U70 ( .A1(n331), .A2(n66), .B1(n328), .B2(n336), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n336) );
  OAI22_X1 U72 ( .A1(n331), .A2(n67), .B1(n328), .B2(n335), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n335) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n368) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module reg_4 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n367), .Z(n329) );
  BUF_X1 U4 ( .A(n367), .Z(n328) );
  BUF_X1 U5 ( .A(n367), .Z(n330) );
  BUF_X1 U6 ( .A(n368), .Z(n331) );
  BUF_X1 U7 ( .A(n368), .Z(n332) );
  BUF_X1 U8 ( .A(n368), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n367) );
  OAI22_X1 U10 ( .A1(n333), .A2(n36), .B1(n330), .B2(n366), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n366) );
  OAI22_X1 U12 ( .A1(n333), .A2(n37), .B1(n330), .B2(n365), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n365) );
  OAI22_X1 U14 ( .A1(n333), .A2(n38), .B1(n330), .B2(n364), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n364) );
  OAI22_X1 U16 ( .A1(n333), .A2(n39), .B1(n330), .B2(n363), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n363) );
  OAI22_X1 U18 ( .A1(n333), .A2(n40), .B1(n330), .B2(n362), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n362) );
  OAI22_X1 U20 ( .A1(n333), .A2(n41), .B1(n330), .B2(n361), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n361) );
  OAI22_X1 U22 ( .A1(n333), .A2(n42), .B1(n330), .B2(n360), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n360) );
  OAI22_X1 U24 ( .A1(n332), .A2(n43), .B1(n330), .B2(n359), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n359) );
  OAI22_X1 U26 ( .A1(n332), .A2(n44), .B1(n329), .B2(n358), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n358) );
  OAI22_X1 U28 ( .A1(n332), .A2(n45), .B1(n329), .B2(n357), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n357) );
  OAI22_X1 U30 ( .A1(n332), .A2(n46), .B1(n329), .B2(n356), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n356) );
  OAI22_X1 U32 ( .A1(n332), .A2(n47), .B1(n329), .B2(n355), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n355) );
  OAI22_X1 U34 ( .A1(n332), .A2(n48), .B1(n329), .B2(n354), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n354) );
  OAI22_X1 U36 ( .A1(n332), .A2(n49), .B1(n329), .B2(n353), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n353) );
  OAI22_X1 U38 ( .A1(n332), .A2(n50), .B1(n329), .B2(n352), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n352) );
  OAI22_X1 U40 ( .A1(n332), .A2(n51), .B1(n329), .B2(n351), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n351) );
  OAI22_X1 U42 ( .A1(n332), .A2(n52), .B1(n329), .B2(n350), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n350) );
  OAI22_X1 U44 ( .A1(n332), .A2(n53), .B1(n329), .B2(n349), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n349) );
  OAI22_X1 U46 ( .A1(n332), .A2(n54), .B1(n329), .B2(n348), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n348) );
  OAI22_X1 U48 ( .A1(n332), .A2(n55), .B1(n329), .B2(n347), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n347) );
  OAI22_X1 U50 ( .A1(n331), .A2(n56), .B1(n328), .B2(n346), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n346) );
  OAI22_X1 U52 ( .A1(n331), .A2(n57), .B1(n328), .B2(n345), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n345) );
  OAI22_X1 U54 ( .A1(n331), .A2(n58), .B1(n328), .B2(n344), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n344) );
  OAI22_X1 U56 ( .A1(n331), .A2(n59), .B1(n328), .B2(n343), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n343) );
  OAI22_X1 U58 ( .A1(n331), .A2(n60), .B1(n328), .B2(n342), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n342) );
  OAI22_X1 U60 ( .A1(n331), .A2(n61), .B1(n328), .B2(n341), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n341) );
  OAI22_X1 U62 ( .A1(n331), .A2(n62), .B1(n328), .B2(n340), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n340) );
  OAI22_X1 U64 ( .A1(n331), .A2(n63), .B1(n328), .B2(n339), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n339) );
  OAI22_X1 U66 ( .A1(n331), .A2(n64), .B1(n328), .B2(n338), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n338) );
  OAI22_X1 U68 ( .A1(n331), .A2(n65), .B1(n328), .B2(n337), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n337) );
  OAI22_X1 U70 ( .A1(n331), .A2(n66), .B1(n328), .B2(n336), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n336) );
  OAI22_X1 U72 ( .A1(n331), .A2(n67), .B1(n328), .B2(n335), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n335) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n368) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module executeUnit_M32_C4 ( clock, reset, en3, Mux1Sel, Mux2Sel, ALUCODE, 
        OUT1RF, OUT2RF, IMMEDIATE, NPCFromDecode, AddressWfromDecode, 
        ALUtoMEMORY, OUT2RFtoMEMORY, AddressWtoMEMORY );
  input [3:0] ALUCODE;
  input [31:0] OUT1RF;
  input [31:0] OUT2RF;
  input [31:0] IMMEDIATE;
  input [31:0] NPCFromDecode;
  input [31:0] AddressWfromDecode;
  output [31:0] ALUtoMEMORY;
  output [31:0] OUT2RFtoMEMORY;
  output [31:0] AddressWtoMEMORY;
  input clock, reset, en3, Mux1Sel, Mux2Sel;

  wire   [31:0] MUX2out;
  wire   [31:0] MUXNPCout;
  wire   [31:0] MUXWITH4out;
  wire   [31:0] ALUout;

  Mux21_4 MUX ( .a(OUT2RF), .b(IMMEDIATE), .sel(Mux2Sel), .y(MUX2out) );
  Mux21_3 MUXNPC ( .a(NPCFromDecode), .b(OUT1RF), .sel(Mux1Sel), .y(MUXNPCout)
         );
  Mux21_2 MUXWITH4 ( .a({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b(MUX2out), .sel(Mux1Sel), .y(MUXWITH4out) );
  ALU_M32_C4 ALUset ( .CODE(ALUCODE), .DATA1(MUXNPCout), .DATA2(MUXWITH4out), 
        .OUTALU(ALUout) );
  reg_6 ALUout_REG ( .clock(clock), .reset(reset), .load(en3), .i(ALUout), .o(
        ALUtoMEMORY) );
  reg_5 RFout2_REG ( .clock(clock), .reset(reset), .load(en3), .i(OUT2RF), .o(
        OUT2RFtoMEMORY) );
  reg_4 AddressW_REG ( .clock(clock), .reset(reset), .load(en3), .i(
        AddressWfromDecode), .o(AddressWtoMEMORY) );
endmodule


module reg_3 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n367), .Z(n329) );
  BUF_X1 U4 ( .A(n367), .Z(n328) );
  BUF_X1 U5 ( .A(n367), .Z(n330) );
  BUF_X1 U6 ( .A(n368), .Z(n331) );
  BUF_X1 U7 ( .A(n368), .Z(n332) );
  BUF_X1 U8 ( .A(n368), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n367) );
  OAI22_X1 U10 ( .A1(n333), .A2(n36), .B1(n330), .B2(n366), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n366) );
  OAI22_X1 U12 ( .A1(n333), .A2(n37), .B1(n330), .B2(n365), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n365) );
  OAI22_X1 U14 ( .A1(n333), .A2(n38), .B1(n330), .B2(n364), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n364) );
  OAI22_X1 U16 ( .A1(n333), .A2(n39), .B1(n330), .B2(n363), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n363) );
  OAI22_X1 U18 ( .A1(n333), .A2(n40), .B1(n330), .B2(n362), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n362) );
  OAI22_X1 U20 ( .A1(n333), .A2(n41), .B1(n330), .B2(n361), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n361) );
  OAI22_X1 U22 ( .A1(n333), .A2(n42), .B1(n330), .B2(n360), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n360) );
  OAI22_X1 U24 ( .A1(n332), .A2(n43), .B1(n330), .B2(n359), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n359) );
  OAI22_X1 U26 ( .A1(n332), .A2(n44), .B1(n329), .B2(n358), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n358) );
  OAI22_X1 U28 ( .A1(n332), .A2(n45), .B1(n329), .B2(n357), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n357) );
  OAI22_X1 U30 ( .A1(n332), .A2(n46), .B1(n329), .B2(n356), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n356) );
  OAI22_X1 U32 ( .A1(n332), .A2(n47), .B1(n329), .B2(n355), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n355) );
  OAI22_X1 U34 ( .A1(n332), .A2(n48), .B1(n329), .B2(n354), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n354) );
  OAI22_X1 U36 ( .A1(n332), .A2(n49), .B1(n329), .B2(n353), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n353) );
  OAI22_X1 U38 ( .A1(n332), .A2(n50), .B1(n329), .B2(n352), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n352) );
  OAI22_X1 U40 ( .A1(n332), .A2(n51), .B1(n329), .B2(n351), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n351) );
  OAI22_X1 U42 ( .A1(n332), .A2(n52), .B1(n329), .B2(n350), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n350) );
  OAI22_X1 U44 ( .A1(n332), .A2(n53), .B1(n329), .B2(n349), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n349) );
  OAI22_X1 U46 ( .A1(n332), .A2(n54), .B1(n329), .B2(n348), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n348) );
  OAI22_X1 U48 ( .A1(n332), .A2(n55), .B1(n329), .B2(n347), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n347) );
  OAI22_X1 U50 ( .A1(n331), .A2(n56), .B1(n328), .B2(n346), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n346) );
  OAI22_X1 U52 ( .A1(n331), .A2(n57), .B1(n328), .B2(n345), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n345) );
  OAI22_X1 U54 ( .A1(n331), .A2(n58), .B1(n328), .B2(n344), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n344) );
  OAI22_X1 U56 ( .A1(n331), .A2(n59), .B1(n328), .B2(n343), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n343) );
  OAI22_X1 U58 ( .A1(n331), .A2(n60), .B1(n328), .B2(n342), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n342) );
  OAI22_X1 U60 ( .A1(n331), .A2(n61), .B1(n328), .B2(n341), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n341) );
  OAI22_X1 U62 ( .A1(n331), .A2(n62), .B1(n328), .B2(n340), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n340) );
  OAI22_X1 U64 ( .A1(n331), .A2(n63), .B1(n328), .B2(n339), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n339) );
  OAI22_X1 U66 ( .A1(n331), .A2(n64), .B1(n328), .B2(n338), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n338) );
  OAI22_X1 U68 ( .A1(n331), .A2(n65), .B1(n328), .B2(n337), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n337) );
  OAI22_X1 U70 ( .A1(n331), .A2(n66), .B1(n328), .B2(n336), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n336) );
  OAI22_X1 U72 ( .A1(n331), .A2(n67), .B1(n328), .B2(n335), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n335) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n368) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module reg_2 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n329) );
  BUF_X1 U4 ( .A(n35), .Z(n328) );
  BUF_X1 U5 ( .A(n35), .Z(n330) );
  BUF_X1 U6 ( .A(n34), .Z(n331) );
  BUF_X1 U7 ( .A(n34), .Z(n332) );
  BUF_X1 U8 ( .A(n34), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n35) );
  OAI22_X1 U10 ( .A1(n333), .A2(n36), .B1(n330), .B2(n335), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n335) );
  OAI22_X1 U12 ( .A1(n333), .A2(n37), .B1(n330), .B2(n336), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n336) );
  OAI22_X1 U14 ( .A1(n333), .A2(n38), .B1(n330), .B2(n337), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n337) );
  OAI22_X1 U16 ( .A1(n333), .A2(n39), .B1(n330), .B2(n338), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n338) );
  OAI22_X1 U18 ( .A1(n333), .A2(n40), .B1(n330), .B2(n339), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n339) );
  OAI22_X1 U20 ( .A1(n333), .A2(n41), .B1(n330), .B2(n340), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n340) );
  OAI22_X1 U22 ( .A1(n333), .A2(n42), .B1(n330), .B2(n341), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n341) );
  OAI22_X1 U24 ( .A1(n332), .A2(n43), .B1(n330), .B2(n342), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n342) );
  OAI22_X1 U26 ( .A1(n332), .A2(n44), .B1(n329), .B2(n343), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n343) );
  OAI22_X1 U28 ( .A1(n332), .A2(n45), .B1(n329), .B2(n344), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n344) );
  OAI22_X1 U30 ( .A1(n332), .A2(n46), .B1(n329), .B2(n345), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n345) );
  OAI22_X1 U32 ( .A1(n332), .A2(n47), .B1(n329), .B2(n346), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n346) );
  OAI22_X1 U34 ( .A1(n332), .A2(n48), .B1(n329), .B2(n347), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n347) );
  OAI22_X1 U36 ( .A1(n332), .A2(n49), .B1(n329), .B2(n348), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n348) );
  OAI22_X1 U38 ( .A1(n332), .A2(n50), .B1(n329), .B2(n349), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n349) );
  OAI22_X1 U40 ( .A1(n332), .A2(n51), .B1(n329), .B2(n350), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n350) );
  OAI22_X1 U42 ( .A1(n332), .A2(n52), .B1(n329), .B2(n351), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n351) );
  OAI22_X1 U44 ( .A1(n332), .A2(n53), .B1(n329), .B2(n352), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n352) );
  OAI22_X1 U46 ( .A1(n332), .A2(n54), .B1(n329), .B2(n353), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n353) );
  OAI22_X1 U48 ( .A1(n332), .A2(n55), .B1(n329), .B2(n354), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n354) );
  OAI22_X1 U50 ( .A1(n331), .A2(n56), .B1(n328), .B2(n355), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n355) );
  OAI22_X1 U52 ( .A1(n331), .A2(n57), .B1(n328), .B2(n356), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n356) );
  OAI22_X1 U54 ( .A1(n331), .A2(n58), .B1(n328), .B2(n357), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n357) );
  OAI22_X1 U56 ( .A1(n331), .A2(n59), .B1(n328), .B2(n358), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n358) );
  OAI22_X1 U58 ( .A1(n331), .A2(n60), .B1(n328), .B2(n359), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n359) );
  OAI22_X1 U60 ( .A1(n331), .A2(n61), .B1(n328), .B2(n360), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n360) );
  OAI22_X1 U62 ( .A1(n331), .A2(n62), .B1(n328), .B2(n361), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n361) );
  OAI22_X1 U64 ( .A1(n331), .A2(n63), .B1(n328), .B2(n362), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n362) );
  OAI22_X1 U66 ( .A1(n331), .A2(n64), .B1(n328), .B2(n363), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n363) );
  OAI22_X1 U68 ( .A1(n331), .A2(n65), .B1(n328), .B2(n364), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n364) );
  OAI22_X1 U70 ( .A1(n331), .A2(n66), .B1(n328), .B2(n365), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n365) );
  OAI22_X1 U72 ( .A1(n331), .A2(n67), .B1(n328), .B2(n366), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n366) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n34) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module reg_1 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n367), .Z(n329) );
  BUF_X1 U4 ( .A(n367), .Z(n328) );
  BUF_X1 U5 ( .A(n367), .Z(n330) );
  BUF_X1 U6 ( .A(n368), .Z(n331) );
  BUF_X1 U7 ( .A(n368), .Z(n332) );
  BUF_X1 U8 ( .A(n368), .Z(n333) );
  NAND2_X1 U9 ( .A1(n334), .A2(n331), .ZN(n367) );
  OAI22_X1 U10 ( .A1(n333), .A2(n36), .B1(n330), .B2(n366), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n366) );
  OAI22_X1 U12 ( .A1(n333), .A2(n37), .B1(n330), .B2(n365), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n365) );
  OAI22_X1 U14 ( .A1(n333), .A2(n38), .B1(n330), .B2(n364), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n364) );
  OAI22_X1 U16 ( .A1(n333), .A2(n39), .B1(n330), .B2(n363), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n363) );
  OAI22_X1 U18 ( .A1(n333), .A2(n40), .B1(n330), .B2(n362), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n362) );
  OAI22_X1 U20 ( .A1(n333), .A2(n41), .B1(n330), .B2(n361), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n361) );
  OAI22_X1 U22 ( .A1(n333), .A2(n42), .B1(n330), .B2(n360), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n360) );
  OAI22_X1 U24 ( .A1(n332), .A2(n43), .B1(n330), .B2(n359), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n359) );
  OAI22_X1 U26 ( .A1(n332), .A2(n44), .B1(n329), .B2(n358), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n358) );
  OAI22_X1 U28 ( .A1(n332), .A2(n45), .B1(n329), .B2(n357), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n357) );
  OAI22_X1 U30 ( .A1(n332), .A2(n46), .B1(n329), .B2(n356), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n356) );
  OAI22_X1 U32 ( .A1(n332), .A2(n47), .B1(n329), .B2(n355), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n355) );
  OAI22_X1 U34 ( .A1(n332), .A2(n48), .B1(n329), .B2(n354), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n354) );
  OAI22_X1 U36 ( .A1(n332), .A2(n49), .B1(n329), .B2(n353), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n353) );
  OAI22_X1 U38 ( .A1(n332), .A2(n50), .B1(n329), .B2(n352), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n352) );
  OAI22_X1 U40 ( .A1(n332), .A2(n51), .B1(n329), .B2(n351), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n351) );
  OAI22_X1 U42 ( .A1(n332), .A2(n52), .B1(n329), .B2(n350), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n350) );
  OAI22_X1 U44 ( .A1(n332), .A2(n53), .B1(n329), .B2(n349), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n349) );
  OAI22_X1 U46 ( .A1(n332), .A2(n54), .B1(n329), .B2(n348), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n348) );
  OAI22_X1 U48 ( .A1(n332), .A2(n55), .B1(n329), .B2(n347), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n347) );
  OAI22_X1 U50 ( .A1(n331), .A2(n56), .B1(n328), .B2(n346), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n346) );
  OAI22_X1 U52 ( .A1(n331), .A2(n57), .B1(n328), .B2(n345), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n345) );
  OAI22_X1 U54 ( .A1(n331), .A2(n58), .B1(n328), .B2(n344), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n344) );
  OAI22_X1 U56 ( .A1(n331), .A2(n59), .B1(n328), .B2(n343), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n343) );
  OAI22_X1 U58 ( .A1(n331), .A2(n60), .B1(n328), .B2(n342), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n342) );
  OAI22_X1 U60 ( .A1(n331), .A2(n61), .B1(n328), .B2(n341), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n341) );
  OAI22_X1 U62 ( .A1(n331), .A2(n62), .B1(n328), .B2(n340), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n340) );
  OAI22_X1 U64 ( .A1(n331), .A2(n63), .B1(n328), .B2(n339), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n339) );
  OAI22_X1 U66 ( .A1(n331), .A2(n64), .B1(n328), .B2(n338), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n338) );
  OAI22_X1 U68 ( .A1(n331), .A2(n65), .B1(n328), .B2(n337), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n337) );
  OAI22_X1 U70 ( .A1(n331), .A2(n66), .B1(n328), .B2(n336), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n336) );
  OAI22_X1 U72 ( .A1(n331), .A2(n67), .B1(n328), .B2(n335), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n335) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n368) );
  INV_X1 U75 ( .A(reset), .ZN(n334) );
endmodule


module memoryUnit ( clock, reset, en4, ALUout, DRAMout, AddressWfromEXECUTE, 
        LOADDATA, ALUtoWBMUX, AddressWtoWB );
  input [31:0] ALUout;
  input [31:0] DRAMout;
  input [31:0] AddressWfromEXECUTE;
  output [31:0] LOADDATA;
  output [31:0] ALUtoWBMUX;
  output [31:0] AddressWtoWB;
  input clock, reset, en4;


  reg_3 LMD_REG ( .clock(clock), .reset(reset), .load(en4), .i(DRAMout), .o(
        LOADDATA) );
  reg_2 ALUout_REG ( .clock(clock), .reset(reset), .load(en4), .i(ALUout), .o(
        ALUtoWBMUX) );
  reg_1 AddressW_REG ( .clock(clock), .reset(reset), .load(en4), .i(
        AddressWfromEXECUTE), .o(AddressWtoWB) );
endmodule


module Mux21_1 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460;

  INV_X1 U1 ( .A(n395), .ZN(n386) );
  BUF_X1 U2 ( .A(n387), .Z(n393) );
  BUF_X1 U3 ( .A(n396), .Z(n391) );
  BUF_X1 U4 ( .A(n396), .Z(n390) );
  BUF_X1 U5 ( .A(n389), .Z(n394) );
  BUF_X1 U6 ( .A(n396), .Z(n392) );
  BUF_X1 U7 ( .A(n396), .Z(n389) );
  BUF_X1 U8 ( .A(n396), .Z(n388) );
  BUF_X1 U9 ( .A(n396), .Z(n387) );
  BUF_X1 U10 ( .A(n396), .Z(n395) );
  INV_X1 U11 ( .A(sel), .ZN(n396) );
  INV_X1 U12 ( .A(n459), .ZN(y[8]) );
  AOI22_X1 U13 ( .A1(a[8]), .A2(n386), .B1(b[8]), .B2(n387), .ZN(n459) );
  INV_X1 U14 ( .A(n453), .ZN(y[31]) );
  AOI22_X1 U15 ( .A1(a[31]), .A2(n386), .B1(b[31]), .B2(n388), .ZN(n453) );
  INV_X1 U16 ( .A(n454), .ZN(y[3]) );
  AOI22_X1 U17 ( .A1(a[3]), .A2(n386), .B1(b[3]), .B2(n388), .ZN(n454) );
  INV_X1 U18 ( .A(n455), .ZN(y[4]) );
  AOI22_X1 U19 ( .A1(a[4]), .A2(n386), .B1(b[4]), .B2(n388), .ZN(n455) );
  INV_X1 U20 ( .A(n456), .ZN(y[5]) );
  AOI22_X1 U21 ( .A1(a[5]), .A2(n386), .B1(b[5]), .B2(n388), .ZN(n456) );
  INV_X1 U22 ( .A(n457), .ZN(y[6]) );
  AOI22_X1 U23 ( .A1(a[6]), .A2(sel), .B1(b[6]), .B2(n387), .ZN(n457) );
  INV_X1 U24 ( .A(n458), .ZN(y[7]) );
  AOI22_X1 U25 ( .A1(a[7]), .A2(sel), .B1(b[7]), .B2(n387), .ZN(n458) );
  INV_X1 U26 ( .A(n460), .ZN(y[9]) );
  AOI22_X1 U27 ( .A1(sel), .A2(a[9]), .B1(b[9]), .B2(n387), .ZN(n460) );
  INV_X1 U28 ( .A(n430), .ZN(y[10]) );
  AOI22_X1 U29 ( .A1(a[10]), .A2(n386), .B1(b[10]), .B2(n394), .ZN(n430) );
  INV_X1 U30 ( .A(n431), .ZN(y[11]) );
  AOI22_X1 U31 ( .A1(a[11]), .A2(n386), .B1(b[11]), .B2(n394), .ZN(n431) );
  INV_X1 U32 ( .A(n432), .ZN(y[12]) );
  AOI22_X1 U33 ( .A1(a[12]), .A2(n386), .B1(b[12]), .B2(n394), .ZN(n432) );
  INV_X1 U34 ( .A(n433), .ZN(y[13]) );
  AOI22_X1 U35 ( .A1(a[13]), .A2(n386), .B1(b[13]), .B2(n393), .ZN(n433) );
  INV_X1 U36 ( .A(n434), .ZN(y[14]) );
  AOI22_X1 U37 ( .A1(a[14]), .A2(n386), .B1(b[14]), .B2(n393), .ZN(n434) );
  INV_X1 U38 ( .A(n435), .ZN(y[15]) );
  AOI22_X1 U39 ( .A1(a[15]), .A2(n386), .B1(b[15]), .B2(n393), .ZN(n435) );
  INV_X1 U40 ( .A(n436), .ZN(y[16]) );
  AOI22_X1 U41 ( .A1(a[16]), .A2(n386), .B1(b[16]), .B2(n393), .ZN(n436) );
  INV_X1 U42 ( .A(n437), .ZN(y[17]) );
  AOI22_X1 U43 ( .A1(a[17]), .A2(n386), .B1(b[17]), .B2(n392), .ZN(n437) );
  INV_X1 U44 ( .A(n438), .ZN(y[18]) );
  AOI22_X1 U45 ( .A1(a[18]), .A2(n386), .B1(b[18]), .B2(n392), .ZN(n438) );
  INV_X1 U46 ( .A(n439), .ZN(y[19]) );
  AOI22_X1 U47 ( .A1(a[19]), .A2(n386), .B1(b[19]), .B2(n392), .ZN(n439) );
  INV_X1 U48 ( .A(n441), .ZN(y[20]) );
  AOI22_X1 U49 ( .A1(a[20]), .A2(sel), .B1(b[20]), .B2(n391), .ZN(n441) );
  INV_X1 U50 ( .A(n442), .ZN(y[21]) );
  AOI22_X1 U51 ( .A1(a[21]), .A2(sel), .B1(b[21]), .B2(n391), .ZN(n442) );
  INV_X1 U52 ( .A(n443), .ZN(y[22]) );
  AOI22_X1 U53 ( .A1(a[22]), .A2(sel), .B1(b[22]), .B2(n391), .ZN(n443) );
  INV_X1 U54 ( .A(n444), .ZN(y[23]) );
  AOI22_X1 U55 ( .A1(a[23]), .A2(sel), .B1(b[23]), .B2(n391), .ZN(n444) );
  INV_X1 U56 ( .A(n445), .ZN(y[24]) );
  AOI22_X1 U57 ( .A1(a[24]), .A2(sel), .B1(b[24]), .B2(n390), .ZN(n445) );
  INV_X1 U58 ( .A(n446), .ZN(y[25]) );
  AOI22_X1 U59 ( .A1(a[25]), .A2(sel), .B1(b[25]), .B2(n390), .ZN(n446) );
  INV_X1 U60 ( .A(n447), .ZN(y[26]) );
  AOI22_X1 U61 ( .A1(a[26]), .A2(sel), .B1(b[26]), .B2(n390), .ZN(n447) );
  INV_X1 U62 ( .A(n448), .ZN(y[27]) );
  AOI22_X1 U63 ( .A1(a[27]), .A2(sel), .B1(b[27]), .B2(n390), .ZN(n448) );
  INV_X1 U64 ( .A(n449), .ZN(y[28]) );
  AOI22_X1 U65 ( .A1(a[28]), .A2(sel), .B1(b[28]), .B2(n389), .ZN(n449) );
  INV_X1 U66 ( .A(n450), .ZN(y[29]) );
  AOI22_X1 U67 ( .A1(a[29]), .A2(sel), .B1(b[29]), .B2(n389), .ZN(n450) );
  INV_X1 U68 ( .A(n452), .ZN(y[30]) );
  AOI22_X1 U69 ( .A1(a[30]), .A2(sel), .B1(b[30]), .B2(n389), .ZN(n452) );
  INV_X1 U70 ( .A(n429), .ZN(y[0]) );
  AOI22_X1 U71 ( .A1(a[0]), .A2(n386), .B1(b[0]), .B2(n394), .ZN(n429) );
  INV_X1 U72 ( .A(n440), .ZN(y[1]) );
  AOI22_X1 U73 ( .A1(a[1]), .A2(n386), .B1(b[1]), .B2(n392), .ZN(n440) );
  INV_X1 U74 ( .A(n451), .ZN(y[2]) );
  AOI22_X1 U75 ( .A1(a[2]), .A2(sel), .B1(b[2]), .B2(n389), .ZN(n451) );
endmodule


module WBUnit ( selwb, ALUin, LOADDATA, AddressWfromMemory, MUXtoRF, 
        AddressWtoDECODE );
  input [31:0] ALUin;
  input [31:0] LOADDATA;
  input [31:0] AddressWfromMemory;
  output [31:0] MUXtoRF;
  output [31:0] AddressWtoDECODE;
  input selwb;

  assign AddressWtoDECODE[31] = AddressWfromMemory[31];
  assign AddressWtoDECODE[30] = AddressWfromMemory[30];
  assign AddressWtoDECODE[29] = AddressWfromMemory[29];
  assign AddressWtoDECODE[28] = AddressWfromMemory[28];
  assign AddressWtoDECODE[27] = AddressWfromMemory[27];
  assign AddressWtoDECODE[26] = AddressWfromMemory[26];
  assign AddressWtoDECODE[25] = AddressWfromMemory[25];
  assign AddressWtoDECODE[24] = AddressWfromMemory[24];
  assign AddressWtoDECODE[23] = AddressWfromMemory[23];
  assign AddressWtoDECODE[22] = AddressWfromMemory[22];
  assign AddressWtoDECODE[21] = AddressWfromMemory[21];
  assign AddressWtoDECODE[20] = AddressWfromMemory[20];
  assign AddressWtoDECODE[19] = AddressWfromMemory[19];
  assign AddressWtoDECODE[18] = AddressWfromMemory[18];
  assign AddressWtoDECODE[17] = AddressWfromMemory[17];
  assign AddressWtoDECODE[16] = AddressWfromMemory[16];
  assign AddressWtoDECODE[15] = AddressWfromMemory[15];
  assign AddressWtoDECODE[14] = AddressWfromMemory[14];
  assign AddressWtoDECODE[13] = AddressWfromMemory[13];
  assign AddressWtoDECODE[12] = AddressWfromMemory[12];
  assign AddressWtoDECODE[11] = AddressWfromMemory[11];
  assign AddressWtoDECODE[10] = AddressWfromMemory[10];
  assign AddressWtoDECODE[9] = AddressWfromMemory[9];
  assign AddressWtoDECODE[8] = AddressWfromMemory[8];
  assign AddressWtoDECODE[7] = AddressWfromMemory[7];
  assign AddressWtoDECODE[6] = AddressWfromMemory[6];
  assign AddressWtoDECODE[5] = AddressWfromMemory[5];
  assign AddressWtoDECODE[4] = AddressWfromMemory[4];
  assign AddressWtoDECODE[3] = AddressWfromMemory[3];
  assign AddressWtoDECODE[2] = AddressWfromMemory[2];
  assign AddressWtoDECODE[1] = AddressWfromMemory[1];
  assign AddressWtoDECODE[0] = AddressWfromMemory[0];

  Mux21_1 wbmux ( .a(LOADDATA), .b(ALUin), .sel(selwb), .y(MUXtoRF) );
endmodule


module dataPath_M32_C4_N5 ( clock, reset, Instruction, en1, en2, SignSelect, 
        RD1, RD2, WR, JMP, BRANCHenable, en3, BranchCondSel, Mux1Sel, Mux2Sel, 
        ALUCODE, RegDestination, en4, DRAMout, selwb, PCtoIM, ALUtoMEMORY, 
        OUT2RFtoMEMORY, InstructionToCU );
  input [31:0] Instruction;
  input [3:0] ALUCODE;
  input [31:0] DRAMout;
  output [31:0] PCtoIM;
  output [31:0] ALUtoMEMORY;
  output [31:0] OUT2RFtoMEMORY;
  output [31:0] InstructionToCU;
  input clock, reset, en1, en2, SignSelect, RD1, RD2, WR, JMP, BRANCHenable,
         en3, BranchCondSel, Mux1Sel, Mux2Sel, RegDestination, en4, selwb;
  wire   BRANCHtoFetch, n1;
  wire   [31:0] NewPC;
  wire   [31:0] NXPC;
  wire   [4:0] AddressfromWB;
  wire   [31:0] MUXtoRF;
  wire   [31:0] OUT1;
  wire   [31:0] OUT2;
  wire   [31:0] OUTIMM;
  wire   [31:0] NPCfromDECODE;
  wire   [31:0] ADDWfromDECODE;
  wire   [31:0] ADDWtoMEMORY;
  wire   [31:0] LOADDATA;
  wire   [31:0] ALUtoWBMUX;
  wire   [31:0] ADDWtoWB;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48;

  fetchUnit FU ( .clock(clock), .reset(n1), .en1(en1), .BranchPC({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, NewPC[9:0]}), 
        .BRANCHfromDECODE(BRANCHtoFetch), .Instruction(Instruction), .PCtoIM(
        PCtoIM), .IRtoDecode(InstructionToCU), .NPCtoDecode(NXPC) );
  DecodeUnit DU ( .clock(clock), .reset(n1), .JMP(JMP), .RegDestination(
        RegDestination), .en2(en2), .SignSelect(SignSelect), .BranchCondSel(
        BranchCondSel), .BRANCHenable(BRANCHenable), .RD1(RD1), .RD2(RD2), 
        .WR(WR), .Instruction(InstructionToCU), .ADD_WR(AddressfromWB), 
        .DATAIN(MUXtoRF), .NPCfromIF(NXPC), .OUT1(OUT1), .OUT2(OUT2), .OUTNPC(
        {SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, NewPC[9:0]}), 
        .OUTIMM(OUTIMM), .NPCtoEX(NPCfromDECODE), .AddressWtoEX(ADDWfromDECODE), .BRANCHtoFetch(BRANCHtoFetch) );
  executeUnit_M32_C4 EU ( .clock(clock), .reset(n1), .en3(en3), .Mux1Sel(
        Mux1Sel), .Mux2Sel(Mux2Sel), .ALUCODE(ALUCODE), .OUT1RF(OUT1), 
        .OUT2RF(OUT2), .IMMEDIATE(OUTIMM), .NPCFromDecode(NPCfromDECODE), 
        .AddressWfromDecode(ADDWfromDECODE), .ALUtoMEMORY(ALUtoMEMORY), 
        .OUT2RFtoMEMORY(OUT2RFtoMEMORY), .AddressWtoMEMORY(ADDWtoMEMORY) );
  memoryUnit MU ( .clock(clock), .reset(n1), .en4(en4), .ALUout(ALUtoMEMORY), 
        .DRAMout(DRAMout), .AddressWfromEXECUTE(ADDWtoMEMORY), .LOADDATA(
        LOADDATA), .ALUtoWBMUX(ALUtoWBMUX), .AddressWtoWB(ADDWtoWB) );
  WBUnit WBU ( .selwb(selwb), .ALUin(ALUtoWBMUX), .LOADDATA(LOADDATA), 
        .AddressWfromMemory(ADDWtoWB), .MUXtoRF(MUXtoRF), .AddressWtoDECODE({
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, AddressfromWB}) );
  BUF_X1 U23 ( .A(reset), .Z(n1) );
endmodule


module DLX_M32_C4_N5 ( Clk, Rst, IRAM_Addr, IRAM_Dout, DRAM_MemoryEnable, 
        DRAM_ReadNotWrite, DRAM_Addr, DRAM_in, DRAM_out );
  output [31:0] IRAM_Addr;
  input [31:0] IRAM_Dout;
  output [4:0] DRAM_Addr;
  output [31:0] DRAM_in;
  input [31:0] DRAM_out;
  input Clk, Rst;
  output DRAM_MemoryEnable, DRAM_ReadNotWrite;
  wire   en2, SignSelect, RD1, RD2, JMP, BranchCondSel, BRANCHenable,
         RegDestination, en3, Mux1Sel, Mux2Sel, en4, selwb, WR;
  wire   [31:0] InstructionToCU;
  wire   [3:0] ALUCODE;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26;

  Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17 CU_I ( .Clk(Clk), .Rst(Rst), .IR_IN(InstructionToCU), .en2(en2), .SignSelect(SignSelect), 
        .RD1(RD1), .RD2(RD2), .JMP(JMP), .BranchCondSel(BranchCondSel), 
        .BRANCHenable(BRANCHenable), .RegDestination(RegDestination), .en3(en3), .Mux1Sel(Mux1Sel), .Mux2Sel(Mux2Sel), .ALUCODE(ALUCODE), .en4(en4), 
        .MemoryEnable(DRAM_MemoryEnable), .ReadNotWrite(DRAM_ReadNotWrite), 
        .selwb(selwb), .WR(WR) );
  dataPath_M32_C4_N5 DP ( .clock(Clk), .reset(Rst), .Instruction(IRAM_Dout), 
        .en1(1'b1), .en2(en2), .SignSelect(SignSelect), .RD1(RD1), .RD2(RD2), 
        .WR(WR), .JMP(JMP), .BRANCHenable(BRANCHenable), .en3(en3), 
        .BranchCondSel(BranchCondSel), .Mux1Sel(Mux1Sel), .Mux2Sel(Mux2Sel), 
        .ALUCODE(ALUCODE), .RegDestination(RegDestination), .en4(en4), 
        .DRAMout(DRAM_out), .selwb(selwb), .PCtoIM(IRAM_Addr), .ALUtoMEMORY({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, DRAM_Addr}), .OUT2RFtoMEMORY(DRAM_in), 
        .InstructionToCU(InstructionToCU) );
endmodule

