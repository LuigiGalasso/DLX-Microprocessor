
module Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17 ( Clk, Rst, 
        IR_IN, en1, en2, SignSelect, RD1, RD2, JMP, BranchCondSel, 
        BRANCHenable, RegDestination, en3, Mux1Sel, Mux2Sel, ALUCODE, en4, 
        MemoryEnable, ReadNotWrite, selwb, WR );
  input [31:0] IR_IN;
  output [3:0] ALUCODE;
  input Clk, Rst;
  output en1, en2, SignSelect, RD1, RD2, JMP, BranchCondSel, BRANCHenable,
         RegDestination, en3, Mux1Sel, Mux2Sel, en4, MemoryEnable,
         ReadNotWrite, selwb, WR;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26, N174,
         N175, N176, N182, N183, N184, N185, n103, n104, n105, n193, n194,
         n195, n275, n276, n277, n278, n279, n280, n281, n282, n283, n358,
         n359, n360, n361, n362, n364, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n363, n365, n366, n367, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n106, n107, n108, n109, n110, n111, n112, n113;
  wire   [7:0] cw2;
  assign en1 = 1'b1;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];

  DFF_X1 \aluOpcode3_reg[3]  ( .D(n105), .CK(Clk), .Q(ALUCODE[3]), .QN(n195)
         );
  DFF_X1 \aluOpcode3_reg[2]  ( .D(n104), .CK(Clk), .Q(ALUCODE[2]), .QN(n194)
         );
  DFF_X1 \aluOpcode3_reg[1]  ( .D(n87), .CK(Clk), .Q(ALUCODE[1]) );
  DLH_X1 \cw2_reg[15]  ( .G(N174), .D(n85), .Q(en2) );
  DLH_X1 \cw2_reg[13]  ( .G(N174), .D(N184), .Q(RD1) );
  DLH_X1 \cw2_reg[12]  ( .G(N174), .D(N183), .Q(RD2) );
  DLH_X1 \cw2_reg[11]  ( .G(N174), .D(N182), .Q(JMP) );
  DLH_X1 \cw2_reg[10]  ( .G(N174), .D(n364), .Q(BranchCondSel) );
  DLH_X1 \cw2_reg[9]  ( .G(N174), .D(n90), .Q(BRANCHenable) );
  DLH_X1 \cw2_reg[8]  ( .G(N174), .D(n88), .Q(RegDestination) );
  DLH_X1 \cw2_reg[7]  ( .G(N174), .D(n85), .Q(cw2[7]) );
  SDFF_X1 \cw3_reg[7]  ( .D(1'b0), .SI(n85), .SE(cw2[7]), .CK(Clk), .Q(en3) );
  DLH_X1 \cw2_reg[6]  ( .G(N174), .D(n91), .Q(cw2[6]) );
  SDFF_X1 \cw3_reg[6]  ( .D(1'b0), .SI(n85), .SE(cw2[6]), .CK(Clk), .Q(Mux1Sel) );
  DLH_X1 \cw2_reg[5]  ( .G(N174), .D(n88), .Q(cw2[5]) );
  DLH_X1 \cw2_reg[4]  ( .G(N174), .D(n85), .Q(cw2[4]) );
  SDFF_X1 \cw3_reg[4]  ( .D(1'b0), .SI(n85), .SE(cw2[4]), .CK(Clk), .QN(n362)
         );
  DLH_X1 \cw2_reg[3]  ( .G(N174), .D(n94), .Q(cw2[3]) );
  SDFF_X1 \cw3_reg[3]  ( .D(1'b0), .SI(n85), .SE(cw2[3]), .CK(Clk), .QN(n361)
         );
  DLH_X1 \cw2_reg[2]  ( .G(N174), .D(N176), .Q(cw2[2]) );
  SDFF_X1 \cw3_reg[2]  ( .D(1'b0), .SI(n85), .SE(cw2[2]), .CK(Clk), .QN(n360)
         );
  DLH_X1 \cw2_reg[1]  ( .G(N174), .D(N176), .Q(cw2[1]) );
  SDFF_X1 \cw3_reg[1]  ( .D(1'b0), .SI(n85), .SE(cw2[1]), .CK(Clk), .QN(n359)
         );
  DLH_X1 \cw2_reg[0]  ( .G(N174), .D(N175), .Q(cw2[0]) );
  SDFF_X1 \cw3_reg[0]  ( .D(1'b0), .SI(n85), .SE(cw2[0]), .CK(Clk), .QN(n358)
         );
  DFF_X1 \cw5_reg[0]  ( .D(n282), .CK(Clk), .Q(WR) );
  DFF_X1 \cw4_reg[4]  ( .D(n281), .CK(Clk), .Q(en4) );
  DFF_X1 \cw4_reg[3]  ( .D(n280), .CK(Clk), .Q(MemoryEnable) );
  DFF_X1 \cw4_reg[2]  ( .D(n279), .CK(Clk), .Q(ReadNotWrite) );
  DFF_X1 \cw4_reg[1]  ( .D(n278), .CK(Clk), .QN(n275) );
  DFF_X1 \cw4_reg[0]  ( .D(n277), .CK(Clk), .QN(n276) );
  OAI33_X1 U296 ( .A1(n111), .A2(n317), .A3(n318), .B1(n319), .B2(n320), .B3(
        n321), .ZN(n316) );
  NAND3_X1 U297 ( .A1(n86), .A2(n320), .A3(n107), .ZN(n331) );
  NAND3_X1 U298 ( .A1(n352), .A2(n349), .A3(n353), .ZN(N174) );
  NAND3_X1 U299 ( .A1(IR_IN_28), .A2(n354), .A3(IR_IN_30), .ZN(n327) );
  NAND3_X1 U300 ( .A1(n365), .A2(n96), .A3(n340), .ZN(n332) );
  NAND3_X1 U301 ( .A1(n366), .A2(n98), .A3(n326), .ZN(n365) );
  NAND3_X1 U302 ( .A1(n340), .A2(n367), .A3(IR_IN_30), .ZN(n330) );
  NAND3_X1 U303 ( .A1(IR_IN_26), .A2(n355), .A3(IR_IN_31), .ZN(n342) );
  SDFF_X1 \cw3_reg[5]  ( .D(1'b0), .SI(n85), .SE(cw2[5]), .CK(Clk), .Q(Mux2Sel) );
  DLH_X1 \cw2_reg[14]  ( .G(N174), .D(N185), .Q(SignSelect) );
  DFF_X1 \cw5_reg[1]  ( .D(n283), .CK(Clk), .Q(selwb) );
  DFF_X1 \aluOpcode3_reg[0]  ( .D(n103), .CK(Clk), .Q(ALUCODE[0]), .QN(n193)
         );
  INV_X1 U210 ( .A(n318), .ZN(n88) );
  INV_X1 U211 ( .A(n321), .ZN(n106) );
  INV_X1 U212 ( .A(n319), .ZN(n86) );
  NAND2_X1 U213 ( .A1(n329), .A2(n318), .ZN(N183) );
  OR2_X1 U214 ( .A1(n88), .A2(N185), .ZN(N184) );
  INV_X1 U215 ( .A(n313), .ZN(n90) );
  INV_X1 U216 ( .A(n329), .ZN(n94) );
  NAND4_X1 U217 ( .A1(n340), .A2(n341), .A3(n99), .A4(n96), .ZN(n343) );
  NAND4_X1 U218 ( .A1(n110), .A2(n109), .A3(n108), .A4(n339), .ZN(n324) );
  NAND2_X1 U219 ( .A1(n348), .A2(n85), .ZN(n318) );
  NAND2_X1 U220 ( .A1(n338), .A2(n110), .ZN(n321) );
  AND3_X1 U221 ( .A1(n351), .A2(n99), .A3(n341), .ZN(n348) );
  AND2_X1 U222 ( .A1(n354), .A2(n96), .ZN(n351) );
  AND2_X1 U223 ( .A1(n354), .A2(n355), .ZN(n346) );
  INV_X1 U224 ( .A(n366), .ZN(n100) );
  INV_X1 U225 ( .A(n340), .ZN(n93) );
  INV_X1 U226 ( .A(n327), .ZN(n92) );
  NAND2_X1 U227 ( .A1(n88), .A2(n112), .ZN(n319) );
  INV_X1 U228 ( .A(n356), .ZN(n98) );
  INV_X1 U229 ( .A(n328), .ZN(n89) );
  NAND2_X1 U230 ( .A1(n111), .A2(n113), .ZN(n320) );
  AOI21_X1 U231 ( .B1(n100), .B2(n351), .A(n95), .ZN(n352) );
  NOR4_X1 U232 ( .A1(Rst), .A2(n348), .A3(n350), .A4(n346), .ZN(n353) );
  AOI21_X1 U233 ( .B1(n85), .B2(n350), .A(n364), .ZN(n313) );
  NAND2_X1 U234 ( .A1(n95), .A2(n85), .ZN(n329) );
  OAI211_X1 U235 ( .C1(Rst), .C2(n349), .A(n329), .B(n313), .ZN(N185) );
  INV_X1 U236 ( .A(n342), .ZN(n95) );
  OAI211_X1 U237 ( .C1(Rst), .C2(n349), .A(n318), .B(n312), .ZN(N175) );
  AND2_X1 U238 ( .A1(n356), .A2(n351), .ZN(n350) );
  AND3_X1 U239 ( .A1(n351), .A2(n85), .A3(n100), .ZN(n364) );
  AND2_X1 U240 ( .A1(n346), .A2(n85), .ZN(N182) );
  INV_X1 U241 ( .A(n312), .ZN(n91) );
  NOR4_X1 U242 ( .A1(IR_IN[9]), .A2(IR_IN[8]), .A3(IR_IN[7]), .A4(IR_IN[6]), 
        .ZN(n339) );
  INV_X1 U243 ( .A(n314), .ZN(n87) );
  AOI221_X1 U244 ( .B1(n315), .B2(n85), .C1(Rst), .C2(ALUCODE[1]), .A(n316), 
        .ZN(n314) );
  OAI221_X1 U245 ( .B1(n98), .B2(n93), .C1(n326), .C2(n327), .A(n89), .ZN(n315) );
  NOR2_X1 U246 ( .A1(n97), .A2(IR_IN_31), .ZN(n340) );
  NOR2_X1 U247 ( .A1(IR_IN_26), .A2(IR_IN_27), .ZN(n341) );
  NOR3_X1 U248 ( .A1(n101), .A2(IR_IN_27), .A3(n99), .ZN(n356) );
  NOR2_X1 U249 ( .A1(n112), .A2(IR_IN[0]), .ZN(n323) );
  OAI221_X1 U250 ( .B1(Rst), .B2(n335), .C1(n193), .C2(n85), .A(n336), .ZN(
        n103) );
  OAI211_X1 U251 ( .C1(n337), .C2(n106), .A(n113), .B(n86), .ZN(n336) );
  AOI221_X1 U252 ( .B1(n340), .B2(n100), .C1(n92), .C2(n341), .A(n328), .ZN(
        n335) );
  AOI21_X1 U253 ( .B1(n324), .B2(n325), .A(n111), .ZN(n337) );
  NAND2_X1 U254 ( .A1(IR_IN_27), .A2(n101), .ZN(n326) );
  NAND4_X1 U255 ( .A1(n342), .A2(n343), .A3(n344), .A4(n345), .ZN(n328) );
  AOI21_X1 U256 ( .B1(IR_IN_26), .B2(n346), .A(n347), .ZN(n345) );
  NAND4_X1 U257 ( .A1(IR_IN[2]), .A2(n323), .A3(n106), .A4(n348), .ZN(n344) );
  NOR4_X1 U258 ( .A1(IR_IN_30), .A2(n99), .A3(n93), .A4(n326), .ZN(n347) );
  NOR2_X1 U259 ( .A1(IR_IN_29), .A2(IR_IN_31), .ZN(n354) );
  AOI22_X1 U260 ( .A1(n322), .A2(IR_IN[0]), .B1(n323), .B2(n102), .ZN(n317) );
  INV_X1 U261 ( .A(n324), .ZN(n102) );
  AOI21_X1 U262 ( .B1(n321), .B2(n325), .A(IR_IN[1]), .ZN(n322) );
  INV_X1 U263 ( .A(IR_IN_28), .ZN(n99) );
  NAND2_X1 U264 ( .A1(IR_IN[3]), .A2(n338), .ZN(n325) );
  NAND2_X1 U265 ( .A1(n341), .A2(IR_IN_28), .ZN(n366) );
  OAI21_X1 U266 ( .B1(IR_IN_27), .B2(n101), .A(n366), .ZN(n367) );
  INV_X1 U267 ( .A(IR_IN_26), .ZN(n101) );
  OAI221_X1 U268 ( .B1(Rst), .B2(n330), .C1(n195), .C2(n85), .A(n331), .ZN(
        n105) );
  INV_X1 U269 ( .A(n325), .ZN(n107) );
  INV_X1 U270 ( .A(IR_IN[1]), .ZN(n112) );
  INV_X1 U271 ( .A(IR_IN_30), .ZN(n96) );
  INV_X1 U272 ( .A(IR_IN[2]), .ZN(n111) );
  INV_X1 U273 ( .A(IR_IN[0]), .ZN(n113) );
  AND4_X1 U274 ( .A1(n108), .A2(n109), .A3(IR_IN[5]), .A4(n339), .ZN(n338) );
  INV_X1 U275 ( .A(IR_IN[3]), .ZN(n110) );
  INV_X1 U276 ( .A(IR_IN_29), .ZN(n97) );
  INV_X1 U277 ( .A(IR_IN[4]), .ZN(n109) );
  INV_X1 U278 ( .A(IR_IN[10]), .ZN(n108) );
  AND3_X1 U279 ( .A1(n99), .A2(n96), .A3(IR_IN_27), .ZN(n355) );
  OAI221_X1 U280 ( .B1(Rst), .B2(n332), .C1(n194), .C2(n85), .A(n333), .ZN(
        n104) );
  OR3_X1 U281 ( .A1(n318), .A2(n334), .A3(n321), .ZN(n333) );
  AOI21_X1 U282 ( .B1(n112), .B2(IR_IN[2]), .A(n323), .ZN(n334) );
  NOR2_X1 U283 ( .A1(Rst), .A2(n358), .ZN(n277) );
  NOR2_X1 U284 ( .A1(Rst), .A2(n359), .ZN(n278) );
  NOR2_X1 U285 ( .A1(Rst), .A2(n360), .ZN(n279) );
  NOR2_X1 U286 ( .A1(Rst), .A2(n361), .ZN(n280) );
  NOR2_X1 U287 ( .A1(Rst), .A2(n362), .ZN(n281) );
  NOR2_X1 U288 ( .A1(Rst), .A2(n276), .ZN(n282) );
  NOR2_X1 U289 ( .A1(Rst), .A2(n275), .ZN(n283) );
  INV_X1 U290 ( .A(Rst), .ZN(n85) );
  NAND2_X1 U291 ( .A1(IR_IN_26), .A2(N182), .ZN(n312) );
  NOR2_X1 U292 ( .A1(IR_IN_29), .A2(n329), .ZN(N176) );
  AND4_X1 U293 ( .A1(n330), .A2(n343), .A3(n332), .A4(n357), .ZN(n349) );
  AOI21_X1 U294 ( .B1(n95), .B2(n97), .A(n363), .ZN(n357) );
  AOI21_X1 U295 ( .B1(IR_IN_27), .B2(n326), .A(n327), .ZN(n363) );
endmodule


module Adder_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;

  wire   [31:1] carry;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module Adder ( A, B, reset, Cin, O, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  input reset, Cin;
  output Cout;
  wire   N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47,
         N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61,
         N62, N63, N64, N65, n7, n8, n9, n10;
  assign Cout = O[31];

  Adder_DW01_add_0 add_1_root_add_26_2 ( .A(A), .B(B), .CI(Cin), .SUM({N65, 
        N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, 
        N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, 
        N36, N35, N34}) );
  BUF_X1 U2 ( .A(n10), .Z(n7) );
  BUF_X1 U3 ( .A(n10), .Z(n8) );
  BUF_X1 U4 ( .A(n10), .Z(n9) );
  AND2_X1 U5 ( .A1(N36), .A2(n8), .ZN(O[2]) );
  AND2_X1 U6 ( .A1(N34), .A2(n7), .ZN(O[0]) );
  AND2_X1 U7 ( .A1(N35), .A2(n7), .ZN(O[1]) );
  AND2_X1 U8 ( .A1(N44), .A2(n7), .ZN(O[10]) );
  AND2_X1 U9 ( .A1(N45), .A2(n7), .ZN(O[11]) );
  AND2_X1 U10 ( .A1(N46), .A2(n7), .ZN(O[12]) );
  AND2_X1 U11 ( .A1(N47), .A2(n7), .ZN(O[13]) );
  AND2_X1 U12 ( .A1(N48), .A2(n7), .ZN(O[14]) );
  AND2_X1 U13 ( .A1(N49), .A2(n7), .ZN(O[15]) );
  AND2_X1 U14 ( .A1(N50), .A2(n7), .ZN(O[16]) );
  AND2_X1 U15 ( .A1(N51), .A2(n7), .ZN(O[17]) );
  AND2_X1 U16 ( .A1(N52), .A2(n7), .ZN(O[18]) );
  AND2_X1 U17 ( .A1(N53), .A2(n7), .ZN(O[19]) );
  AND2_X1 U18 ( .A1(N54), .A2(n8), .ZN(O[20]) );
  AND2_X1 U19 ( .A1(N55), .A2(n8), .ZN(O[21]) );
  AND2_X1 U20 ( .A1(N56), .A2(n8), .ZN(O[22]) );
  AND2_X1 U21 ( .A1(N57), .A2(n8), .ZN(O[23]) );
  AND2_X1 U22 ( .A1(N58), .A2(n8), .ZN(O[24]) );
  AND2_X1 U23 ( .A1(N59), .A2(n8), .ZN(O[25]) );
  AND2_X1 U24 ( .A1(N60), .A2(n8), .ZN(O[26]) );
  AND2_X1 U25 ( .A1(N61), .A2(n8), .ZN(O[27]) );
  AND2_X1 U26 ( .A1(N62), .A2(n8), .ZN(O[28]) );
  AND2_X1 U27 ( .A1(N63), .A2(n8), .ZN(O[29]) );
  AND2_X1 U28 ( .A1(N64), .A2(n8), .ZN(O[30]) );
  AND2_X1 U29 ( .A1(N41), .A2(n9), .ZN(O[7]) );
  AND2_X1 U30 ( .A1(N40), .A2(n9), .ZN(O[6]) );
  AND2_X1 U31 ( .A1(N39), .A2(n9), .ZN(O[5]) );
  AND2_X1 U32 ( .A1(N43), .A2(n9), .ZN(O[9]) );
  AND2_X1 U33 ( .A1(N42), .A2(n9), .ZN(O[8]) );
  AND2_X1 U34 ( .A1(N37), .A2(n9), .ZN(O[3]) );
  AND2_X1 U35 ( .A1(N38), .A2(n9), .ZN(O[4]) );
  INV_X1 U36 ( .A(reset), .ZN(n10) );
  AND2_X1 U37 ( .A1(N65), .A2(n9), .ZN(O[31]) );
endmodule


module Mux21_0 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158;

  INV_X1 U1 ( .A(n157), .ZN(n145) );
  CLKBUF_X1 U2 ( .A(n158), .Z(n156) );
  CLKBUF_X1 U3 ( .A(n158), .Z(n155) );
  INV_X1 U4 ( .A(n157), .ZN(n148) );
  INV_X1 U5 ( .A(n157), .ZN(n147) );
  BUF_X1 U6 ( .A(n158), .Z(n157) );
  BUF_X1 U7 ( .A(n158), .Z(n154) );
  BUF_X1 U8 ( .A(n154), .Z(n149) );
  BUF_X1 U9 ( .A(n158), .Z(n153) );
  BUF_X1 U10 ( .A(n158), .Z(n152) );
  BUF_X1 U11 ( .A(n153), .Z(n151) );
  BUF_X1 U12 ( .A(n152), .Z(n150) );
  INV_X1 U13 ( .A(n146), .ZN(n158) );
  BUF_X1 U14 ( .A(sel), .Z(n146) );
  INV_X1 U15 ( .A(n43), .ZN(y[2]) );
  AOI22_X1 U16 ( .A1(a[2]), .A2(n148), .B1(b[2]), .B2(n151), .ZN(n43) );
  INV_X1 U17 ( .A(n64), .ZN(y[10]) );
  AOI22_X1 U18 ( .A1(a[10]), .A2(n148), .B1(b[10]), .B2(n156), .ZN(n64) );
  INV_X1 U19 ( .A(n63), .ZN(y[11]) );
  AOI22_X1 U20 ( .A1(a[11]), .A2(n147), .B1(b[11]), .B2(n156), .ZN(n63) );
  INV_X1 U21 ( .A(n62), .ZN(y[12]) );
  AOI22_X1 U22 ( .A1(a[12]), .A2(n145), .B1(b[12]), .B2(n156), .ZN(n62) );
  INV_X1 U23 ( .A(n61), .ZN(y[13]) );
  AOI22_X1 U24 ( .A1(a[13]), .A2(n147), .B1(b[13]), .B2(n155), .ZN(n61) );
  INV_X1 U25 ( .A(n60), .ZN(y[14]) );
  AOI22_X1 U26 ( .A1(a[14]), .A2(n145), .B1(b[14]), .B2(n155), .ZN(n60) );
  INV_X1 U27 ( .A(n59), .ZN(y[15]) );
  AOI22_X1 U28 ( .A1(a[15]), .A2(n147), .B1(b[15]), .B2(n155), .ZN(n59) );
  INV_X1 U29 ( .A(n58), .ZN(y[16]) );
  AOI22_X1 U30 ( .A1(a[16]), .A2(n145), .B1(b[16]), .B2(n155), .ZN(n58) );
  INV_X1 U31 ( .A(n57), .ZN(y[17]) );
  AOI22_X1 U32 ( .A1(a[17]), .A2(n147), .B1(b[17]), .B2(n154), .ZN(n57) );
  INV_X1 U33 ( .A(n65), .ZN(y[0]) );
  AOI22_X1 U34 ( .A1(a[0]), .A2(n148), .B1(b[0]), .B2(n156), .ZN(n65) );
  INV_X1 U35 ( .A(n54), .ZN(y[1]) );
  AOI22_X1 U36 ( .A1(a[1]), .A2(n148), .B1(b[1]), .B2(n154), .ZN(n54) );
  INV_X1 U37 ( .A(n36), .ZN(y[7]) );
  AOI22_X1 U38 ( .A1(a[7]), .A2(n145), .B1(b[7]), .B2(n149), .ZN(n36) );
  INV_X1 U39 ( .A(n37), .ZN(y[6]) );
  AOI22_X1 U40 ( .A1(a[6]), .A2(n147), .B1(b[6]), .B2(n149), .ZN(n37) );
  INV_X1 U41 ( .A(n38), .ZN(y[5]) );
  AOI22_X1 U42 ( .A1(a[5]), .A2(n145), .B1(b[5]), .B2(n150), .ZN(n38) );
  INV_X1 U43 ( .A(n35), .ZN(y[8]) );
  AOI22_X1 U44 ( .A1(a[8]), .A2(n147), .B1(b[8]), .B2(n149), .ZN(n35) );
  INV_X1 U45 ( .A(n40), .ZN(y[3]) );
  AOI22_X1 U46 ( .A1(a[3]), .A2(n145), .B1(b[3]), .B2(n150), .ZN(n40) );
  INV_X1 U47 ( .A(n34), .ZN(y[9]) );
  AOI22_X1 U48 ( .A1(n147), .A2(a[9]), .B1(b[9]), .B2(n149), .ZN(n34) );
  INV_X1 U49 ( .A(n39), .ZN(y[4]) );
  INV_X1 U50 ( .A(n56), .ZN(y[18]) );
  AOI22_X1 U51 ( .A1(a[18]), .A2(n148), .B1(b[18]), .B2(n154), .ZN(n56) );
  INV_X1 U52 ( .A(n55), .ZN(y[19]) );
  AOI22_X1 U53 ( .A1(a[19]), .A2(n148), .B1(b[19]), .B2(n154), .ZN(n55) );
  INV_X1 U54 ( .A(n53), .ZN(y[20]) );
  AOI22_X1 U55 ( .A1(a[20]), .A2(n148), .B1(b[20]), .B2(n153), .ZN(n53) );
  INV_X1 U56 ( .A(n52), .ZN(y[21]) );
  AOI22_X1 U57 ( .A1(a[21]), .A2(n145), .B1(b[21]), .B2(n153), .ZN(n52) );
  INV_X1 U58 ( .A(n51), .ZN(y[22]) );
  AOI22_X1 U59 ( .A1(a[22]), .A2(n148), .B1(b[22]), .B2(n153), .ZN(n51) );
  INV_X1 U60 ( .A(n50), .ZN(y[23]) );
  AOI22_X1 U61 ( .A1(a[23]), .A2(n147), .B1(b[23]), .B2(n153), .ZN(n50) );
  INV_X1 U62 ( .A(n49), .ZN(y[24]) );
  AOI22_X1 U63 ( .A1(a[24]), .A2(n148), .B1(b[24]), .B2(n152), .ZN(n49) );
  INV_X1 U64 ( .A(n48), .ZN(y[25]) );
  AOI22_X1 U65 ( .A1(a[25]), .A2(n145), .B1(b[25]), .B2(n152), .ZN(n48) );
  INV_X1 U66 ( .A(n47), .ZN(y[26]) );
  AOI22_X1 U67 ( .A1(a[26]), .A2(n145), .B1(b[26]), .B2(n152), .ZN(n47) );
  INV_X1 U68 ( .A(n46), .ZN(y[27]) );
  AOI22_X1 U69 ( .A1(a[27]), .A2(n147), .B1(b[27]), .B2(n152), .ZN(n46) );
  INV_X1 U70 ( .A(n45), .ZN(y[28]) );
  AOI22_X1 U71 ( .A1(a[28]), .A2(n148), .B1(b[28]), .B2(n151), .ZN(n45) );
  INV_X1 U72 ( .A(n44), .ZN(y[29]) );
  AOI22_X1 U73 ( .A1(a[29]), .A2(n145), .B1(b[29]), .B2(n151), .ZN(n44) );
  INV_X1 U74 ( .A(n42), .ZN(y[30]) );
  AOI22_X1 U75 ( .A1(a[30]), .A2(n148), .B1(b[30]), .B2(n151), .ZN(n42) );
  INV_X1 U76 ( .A(n41), .ZN(y[31]) );
  AOI22_X1 U77 ( .A1(a[31]), .A2(n147), .B1(b[31]), .B2(n150), .ZN(n41) );
  AOI22_X1 U78 ( .A1(a[4]), .A2(n145), .B1(b[4]), .B2(n150), .ZN(n39) );
endmodule


module IR ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n31, n32, n33, n34, n35, n97, n98, n99, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n64) );
  DFF_X1 \temp_reg[30]  ( .D(n67), .CK(clock), .Q(o[30]), .QN(n97) );
  DFF_X1 \temp_reg[29]  ( .D(n69), .CK(clock), .Q(o[29]), .QN(n63) );
  DFF_X1 \temp_reg[28]  ( .D(n66), .CK(clock), .Q(o[28]), .QN(n98) );
  DFF_X1 \temp_reg[27]  ( .D(n70), .CK(clock), .Q(o[27]), .QN(n62) );
  DFF_X1 \temp_reg[26]  ( .D(n65), .CK(clock), .Q(o[26]), .QN(n99) );
  DFF_X1 \temp_reg[24]  ( .D(n72), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n73), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n74), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n75), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n76), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n77), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n78), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n79), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n80), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n81), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n82), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n83), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n84), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n85), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n86), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n87), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n88), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n89), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n90), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n91), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n92), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n93), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n94), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n95), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n96), .CK(clock), .Q(o[0]), .QN(n36) );
  DFF_X1 \temp_reg[25]  ( .D(n71), .CK(clock), .Q(o[25]), .QN(n61) );
  BUF_X1 U3 ( .A(n32), .Z(n171) );
  BUF_X1 U4 ( .A(n32), .Z(n172) );
  BUF_X1 U5 ( .A(n32), .Z(n173) );
  INV_X1 U6 ( .A(reset), .ZN(n177) );
  NAND2_X1 U7 ( .A1(n177), .A2(n174), .ZN(n32) );
  BUF_X1 U8 ( .A(n31), .Z(n174) );
  BUF_X1 U9 ( .A(n31), .Z(n175) );
  BUF_X1 U10 ( .A(n31), .Z(n176) );
  OAI22_X1 U11 ( .A1(n175), .A2(n36), .B1(n171), .B2(n206), .ZN(n96) );
  INV_X1 U12 ( .A(i[0]), .ZN(n206) );
  OAI22_X1 U13 ( .A1(n174), .A2(n37), .B1(n171), .B2(n205), .ZN(n95) );
  INV_X1 U14 ( .A(i[1]), .ZN(n205) );
  OAI22_X1 U15 ( .A1(n174), .A2(n38), .B1(n171), .B2(n204), .ZN(n94) );
  INV_X1 U16 ( .A(i[2]), .ZN(n204) );
  OAI22_X1 U17 ( .A1(n174), .A2(n39), .B1(n171), .B2(n203), .ZN(n93) );
  INV_X1 U18 ( .A(i[3]), .ZN(n203) );
  OAI22_X1 U19 ( .A1(n174), .A2(n40), .B1(n171), .B2(n202), .ZN(n92) );
  INV_X1 U20 ( .A(i[4]), .ZN(n202) );
  OAI22_X1 U21 ( .A1(n174), .A2(n41), .B1(n171), .B2(n201), .ZN(n91) );
  INV_X1 U22 ( .A(i[5]), .ZN(n201) );
  OAI22_X1 U23 ( .A1(n174), .A2(n42), .B1(n171), .B2(n200), .ZN(n90) );
  INV_X1 U24 ( .A(i[6]), .ZN(n200) );
  OAI22_X1 U25 ( .A1(n174), .A2(n43), .B1(n171), .B2(n199), .ZN(n89) );
  INV_X1 U26 ( .A(i[7]), .ZN(n199) );
  OAI22_X1 U27 ( .A1(n174), .A2(n44), .B1(n171), .B2(n198), .ZN(n88) );
  INV_X1 U28 ( .A(i[8]), .ZN(n198) );
  OAI22_X1 U29 ( .A1(n174), .A2(n45), .B1(n171), .B2(n197), .ZN(n87) );
  INV_X1 U30 ( .A(i[9]), .ZN(n197) );
  OAI22_X1 U31 ( .A1(n175), .A2(n46), .B1(n171), .B2(n196), .ZN(n86) );
  INV_X1 U32 ( .A(i[10]), .ZN(n196) );
  OAI22_X1 U33 ( .A1(n175), .A2(n47), .B1(n171), .B2(n195), .ZN(n85) );
  INV_X1 U34 ( .A(i[11]), .ZN(n195) );
  OAI22_X1 U35 ( .A1(n175), .A2(n48), .B1(n172), .B2(n194), .ZN(n84) );
  INV_X1 U36 ( .A(i[12]), .ZN(n194) );
  OAI22_X1 U37 ( .A1(n175), .A2(n49), .B1(n172), .B2(n193), .ZN(n83) );
  INV_X1 U38 ( .A(i[13]), .ZN(n193) );
  OAI22_X1 U39 ( .A1(n175), .A2(n50), .B1(n172), .B2(n192), .ZN(n82) );
  INV_X1 U40 ( .A(i[14]), .ZN(n192) );
  OAI22_X1 U41 ( .A1(n175), .A2(n51), .B1(n172), .B2(n191), .ZN(n81) );
  INV_X1 U42 ( .A(i[15]), .ZN(n191) );
  OAI22_X1 U43 ( .A1(n175), .A2(n52), .B1(n172), .B2(n190), .ZN(n80) );
  INV_X1 U44 ( .A(i[16]), .ZN(n190) );
  OAI22_X1 U45 ( .A1(n175), .A2(n53), .B1(n172), .B2(n189), .ZN(n79) );
  INV_X1 U46 ( .A(i[17]), .ZN(n189) );
  OAI22_X1 U47 ( .A1(n175), .A2(n54), .B1(n172), .B2(n188), .ZN(n78) );
  INV_X1 U48 ( .A(i[18]), .ZN(n188) );
  OAI22_X1 U49 ( .A1(n175), .A2(n55), .B1(n172), .B2(n187), .ZN(n77) );
  INV_X1 U50 ( .A(i[19]), .ZN(n187) );
  OAI22_X1 U51 ( .A1(n175), .A2(n56), .B1(n172), .B2(n186), .ZN(n76) );
  INV_X1 U52 ( .A(i[20]), .ZN(n186) );
  OAI22_X1 U53 ( .A1(n175), .A2(n57), .B1(n172), .B2(n185), .ZN(n75) );
  INV_X1 U54 ( .A(i[21]), .ZN(n185) );
  OAI22_X1 U55 ( .A1(n176), .A2(n58), .B1(n172), .B2(n184), .ZN(n74) );
  INV_X1 U56 ( .A(i[22]), .ZN(n184) );
  OAI22_X1 U57 ( .A1(n176), .A2(n59), .B1(n172), .B2(n183), .ZN(n73) );
  INV_X1 U58 ( .A(i[23]), .ZN(n183) );
  OAI22_X1 U59 ( .A1(n176), .A2(n61), .B1(n173), .B2(n181), .ZN(n71) );
  INV_X1 U60 ( .A(i[25]), .ZN(n181) );
  OAI22_X1 U61 ( .A1(n176), .A2(n60), .B1(n173), .B2(n182), .ZN(n72) );
  INV_X1 U62 ( .A(i[24]), .ZN(n182) );
  OAI22_X1 U63 ( .A1(n176), .A2(n62), .B1(n173), .B2(n180), .ZN(n70) );
  INV_X1 U64 ( .A(i[27]), .ZN(n180) );
  OAI22_X1 U65 ( .A1(n176), .A2(n63), .B1(n173), .B2(n179), .ZN(n69) );
  INV_X1 U66 ( .A(i[29]), .ZN(n179) );
  OAI22_X1 U67 ( .A1(n176), .A2(n64), .B1(n173), .B2(n178), .ZN(n68) );
  INV_X1 U68 ( .A(i[31]), .ZN(n178) );
  OAI211_X1 U69 ( .C1(n176), .C2(n99), .A(n35), .B(n177), .ZN(n65) );
  NAND2_X1 U70 ( .A1(i[26]), .A2(n174), .ZN(n35) );
  OAI211_X1 U71 ( .C1(n176), .C2(n98), .A(n34), .B(n177), .ZN(n66) );
  NAND2_X1 U72 ( .A1(i[28]), .A2(n174), .ZN(n34) );
  OAI211_X1 U73 ( .C1(n176), .C2(n97), .A(n33), .B(n177), .ZN(n67) );
  NAND2_X1 U74 ( .A1(i[30]), .A2(n174), .ZN(n33) );
  OR2_X1 U75 ( .A1(reset), .A2(load), .ZN(n31) );
endmodule


module reg_0 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212;

  DFF_X1 \temp_reg[31]  ( .D(n78), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n79), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n80), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n81), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n82), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n83), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n84), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n85), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n86), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n87), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n88), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n89), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n90), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n91), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n92), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n93), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n94), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n95), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n96), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n97), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n98), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n99), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[3]  ( .D(n74), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[1]  ( .D(n76), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[8]  ( .D(n69), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[9]  ( .D(n68), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[0]  ( .D(n77), .CK(clock), .Q(o[0]), .QN(n36) );
  DFF_X1 \temp_reg[5]  ( .D(n72), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[6]  ( .D(n71), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[7]  ( .D(n70), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[4]  ( .D(n73), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[2]  ( .D(n75), .CK(clock), .Q(o[2]), .QN(n38) );
  BUF_X1 U3 ( .A(n35), .Z(n175) );
  BUF_X1 U4 ( .A(n35), .Z(n174) );
  BUF_X1 U5 ( .A(n35), .Z(n176) );
  BUF_X1 U6 ( .A(n34), .Z(n178) );
  BUF_X1 U7 ( .A(n34), .Z(n177) );
  BUF_X1 U8 ( .A(n34), .Z(n179) );
  NAND2_X1 U9 ( .A1(n180), .A2(n177), .ZN(n35) );
  INV_X1 U10 ( .A(i[2]), .ZN(n190) );
  OAI22_X1 U11 ( .A1(n179), .A2(n46), .B1(n176), .B2(n211), .ZN(n99) );
  INV_X1 U12 ( .A(i[10]), .ZN(n211) );
  OAI22_X1 U13 ( .A1(n179), .A2(n47), .B1(n176), .B2(n210), .ZN(n98) );
  INV_X1 U14 ( .A(i[11]), .ZN(n210) );
  OAI22_X1 U15 ( .A1(n179), .A2(n48), .B1(n176), .B2(n209), .ZN(n97) );
  INV_X1 U16 ( .A(i[12]), .ZN(n209) );
  OAI22_X1 U17 ( .A1(n179), .A2(n49), .B1(n176), .B2(n208), .ZN(n96) );
  INV_X1 U18 ( .A(i[13]), .ZN(n208) );
  OAI22_X1 U19 ( .A1(n179), .A2(n50), .B1(n176), .B2(n207), .ZN(n95) );
  INV_X1 U20 ( .A(i[14]), .ZN(n207) );
  OAI22_X1 U21 ( .A1(n179), .A2(n51), .B1(n176), .B2(n206), .ZN(n94) );
  INV_X1 U22 ( .A(i[15]), .ZN(n206) );
  OAI22_X1 U23 ( .A1(n179), .A2(n52), .B1(n176), .B2(n205), .ZN(n93) );
  INV_X1 U24 ( .A(i[16]), .ZN(n205) );
  OAI22_X1 U25 ( .A1(n178), .A2(n53), .B1(n176), .B2(n204), .ZN(n92) );
  INV_X1 U26 ( .A(i[17]), .ZN(n204) );
  OAI22_X1 U27 ( .A1(n177), .A2(n36), .B1(n174), .B2(n212), .ZN(n77) );
  INV_X1 U28 ( .A(i[0]), .ZN(n212) );
  OAI22_X1 U29 ( .A1(n177), .A2(n37), .B1(n174), .B2(n201), .ZN(n76) );
  INV_X1 U30 ( .A(i[1]), .ZN(n201) );
  OAI22_X1 U31 ( .A1(n177), .A2(n43), .B1(n174), .B2(n183), .ZN(n70) );
  INV_X1 U32 ( .A(i[7]), .ZN(n183) );
  OAI22_X1 U33 ( .A1(n177), .A2(n42), .B1(n174), .B2(n184), .ZN(n71) );
  INV_X1 U34 ( .A(i[6]), .ZN(n184) );
  OAI22_X1 U35 ( .A1(n177), .A2(n41), .B1(n174), .B2(n185), .ZN(n72) );
  INV_X1 U36 ( .A(i[5]), .ZN(n185) );
  OAI22_X1 U37 ( .A1(n177), .A2(n44), .B1(n174), .B2(n182), .ZN(n69) );
  INV_X1 U38 ( .A(i[8]), .ZN(n182) );
  OAI22_X1 U39 ( .A1(n177), .A2(n39), .B1(n174), .B2(n187), .ZN(n74) );
  INV_X1 U40 ( .A(i[3]), .ZN(n187) );
  OAI22_X1 U41 ( .A1(n177), .A2(n45), .B1(n174), .B2(n181), .ZN(n68) );
  INV_X1 U42 ( .A(i[9]), .ZN(n181) );
  OAI22_X1 U43 ( .A1(n177), .A2(n40), .B1(n174), .B2(n186), .ZN(n73) );
  INV_X1 U44 ( .A(i[4]), .ZN(n186) );
  OAI22_X1 U45 ( .A1(n178), .A2(n54), .B1(n175), .B2(n203), .ZN(n91) );
  INV_X1 U46 ( .A(i[18]), .ZN(n203) );
  OAI22_X1 U47 ( .A1(n178), .A2(n55), .B1(n175), .B2(n202), .ZN(n90) );
  INV_X1 U48 ( .A(i[19]), .ZN(n202) );
  OAI22_X1 U49 ( .A1(n178), .A2(n56), .B1(n175), .B2(n200), .ZN(n89) );
  INV_X1 U50 ( .A(i[20]), .ZN(n200) );
  OAI22_X1 U51 ( .A1(n178), .A2(n57), .B1(n175), .B2(n199), .ZN(n88) );
  INV_X1 U52 ( .A(i[21]), .ZN(n199) );
  OAI22_X1 U53 ( .A1(n178), .A2(n58), .B1(n175), .B2(n198), .ZN(n87) );
  INV_X1 U54 ( .A(i[22]), .ZN(n198) );
  OAI22_X1 U55 ( .A1(n178), .A2(n59), .B1(n175), .B2(n197), .ZN(n86) );
  INV_X1 U56 ( .A(i[23]), .ZN(n197) );
  OAI22_X1 U57 ( .A1(n178), .A2(n60), .B1(n175), .B2(n196), .ZN(n85) );
  INV_X1 U58 ( .A(i[24]), .ZN(n196) );
  OAI22_X1 U59 ( .A1(n178), .A2(n61), .B1(n175), .B2(n195), .ZN(n84) );
  INV_X1 U60 ( .A(i[25]), .ZN(n195) );
  OAI22_X1 U61 ( .A1(n178), .A2(n62), .B1(n175), .B2(n194), .ZN(n83) );
  INV_X1 U62 ( .A(i[26]), .ZN(n194) );
  OAI22_X1 U63 ( .A1(n178), .A2(n63), .B1(n175), .B2(n193), .ZN(n82) );
  INV_X1 U64 ( .A(i[27]), .ZN(n193) );
  OAI22_X1 U65 ( .A1(n178), .A2(n64), .B1(n175), .B2(n192), .ZN(n81) );
  INV_X1 U66 ( .A(i[28]), .ZN(n192) );
  OAI22_X1 U67 ( .A1(n178), .A2(n65), .B1(n175), .B2(n191), .ZN(n80) );
  INV_X1 U68 ( .A(i[29]), .ZN(n191) );
  OAI22_X1 U69 ( .A1(n177), .A2(n66), .B1(n174), .B2(n189), .ZN(n79) );
  INV_X1 U70 ( .A(i[30]), .ZN(n189) );
  OAI22_X1 U71 ( .A1(n177), .A2(n67), .B1(n174), .B2(n188), .ZN(n78) );
  INV_X1 U72 ( .A(i[31]), .ZN(n188) );
  OR2_X1 U73 ( .A1(load), .A2(reset), .ZN(n34) );
  OAI22_X1 U74 ( .A1(n177), .A2(n38), .B1(n174), .B2(n190), .ZN(n75) );
  INV_X1 U75 ( .A(reset), .ZN(n180) );
endmodule


module reg_12 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n177) );
  BUF_X1 U4 ( .A(n35), .Z(n176) );
  BUF_X1 U5 ( .A(n35), .Z(n178) );
  BUF_X1 U6 ( .A(n34), .Z(n179) );
  BUF_X1 U7 ( .A(n34), .Z(n180) );
  BUF_X1 U8 ( .A(n34), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n35) );
  OAI22_X1 U10 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U12 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n213) );
  OAI22_X1 U14 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U16 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U18 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U20 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U22 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U24 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U26 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U28 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n205) );
  OAI22_X1 U30 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U32 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U34 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U36 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U38 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U40 ( .A1(n180), .A2(n51), .B1(n177), .B2(n199), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n199) );
  OAI22_X1 U42 ( .A1(n180), .A2(n52), .B1(n177), .B2(n198), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n198) );
  OAI22_X1 U44 ( .A1(n180), .A2(n53), .B1(n177), .B2(n197), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n197) );
  OAI22_X1 U46 ( .A1(n180), .A2(n54), .B1(n177), .B2(n196), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n196) );
  OAI22_X1 U48 ( .A1(n180), .A2(n55), .B1(n177), .B2(n195), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n195) );
  OAI22_X1 U50 ( .A1(n179), .A2(n56), .B1(n176), .B2(n194), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n194) );
  OAI22_X1 U52 ( .A1(n179), .A2(n57), .B1(n176), .B2(n193), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n193) );
  OAI22_X1 U54 ( .A1(n179), .A2(n58), .B1(n176), .B2(n192), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n192) );
  OAI22_X1 U56 ( .A1(n179), .A2(n59), .B1(n176), .B2(n191), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n191) );
  OAI22_X1 U58 ( .A1(n179), .A2(n60), .B1(n176), .B2(n190), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n190) );
  OAI22_X1 U60 ( .A1(n179), .A2(n61), .B1(n176), .B2(n189), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n189) );
  OAI22_X1 U62 ( .A1(n179), .A2(n62), .B1(n176), .B2(n188), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n188) );
  OAI22_X1 U64 ( .A1(n179), .A2(n63), .B1(n176), .B2(n187), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n187) );
  OAI22_X1 U66 ( .A1(n179), .A2(n64), .B1(n176), .B2(n186), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n186) );
  OAI22_X1 U68 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U70 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U72 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n183) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n34) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module fetchUnit ( clock, reset, en1, BranchPC, BRANCHfromDECODE, Instruction, 
        PCtoIM, IRtoDecode, NPCtoDecode );
  input [31:0] BranchPC;
  input [31:0] Instruction;
  output [31:0] PCtoIM;
  output [31:0] IRtoDecode;
  output [31:0] NPCtoDecode;
  input clock, reset, en1, BRANCHfromDECODE;
  wire   LOAD;
  wire   [31:0] AddertoMux;
  wire   [31:0] MuxtoPc;

  Adder nxpc ( .A(PCtoIM), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .reset(reset), .Cin(1'b0), .O(AddertoMux) );
  Mux21_0 pcmux ( .a(BranchPC), .b(AddertoMux), .sel(BRANCHfromDECODE), .y(
        MuxtoPc) );
  IR InstrReg ( .clock(clock), .reset(LOAD), .load(en1), .i(Instruction), .o(
        IRtoDecode) );
  reg_0 PC ( .clock(clock), .reset(reset), .load(en1), .i(MuxtoPc), .o(PCtoIM)
         );
  reg_12 NPC ( .clock(clock), .reset(reset), .load(en1), .i(AddertoMux), .o(
        NPCtoDecode) );
  OR2_X1 U2 ( .A1(BRANCHfromDECODE), .A2(reset), .ZN(LOAD) );
endmodule


module Mux41 ( a, b, c, d, sel, y );
  input [31:0] a;
  input [31:0] b;
  input [31:0] c;
  input [31:0] d;
  input [1:0] sel;
  output [31:0] y;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166;

  BUF_X1 U1 ( .A(n6), .Z(n157) );
  BUF_X1 U2 ( .A(n6), .Z(n158) );
  BUF_X1 U3 ( .A(n4), .Z(n163) );
  BUF_X1 U4 ( .A(n4), .Z(n164) );
  BUF_X1 U5 ( .A(n7), .Z(n154) );
  BUF_X1 U6 ( .A(n7), .Z(n155) );
  BUF_X1 U7 ( .A(n5), .Z(n160) );
  BUF_X1 U8 ( .A(n5), .Z(n161) );
  BUF_X1 U9 ( .A(n6), .Z(n159) );
  BUF_X1 U10 ( .A(n4), .Z(n165) );
  BUF_X1 U11 ( .A(n7), .Z(n156) );
  BUF_X1 U12 ( .A(n5), .Z(n162) );
  AOI22_X1 U13 ( .A1(a[4]), .A2(n159), .B1(b[4]), .B2(n156), .ZN(n16) );
  NAND2_X1 U14 ( .A1(n68), .A2(n69), .ZN(y[0]) );
  AOI22_X1 U15 ( .A1(c[0]), .A2(n163), .B1(d[0]), .B2(n160), .ZN(n69) );
  NAND2_X1 U16 ( .A1(n16), .A2(n17), .ZN(y[4]) );
  AOI22_X1 U17 ( .A1(c[4]), .A2(n165), .B1(d[4]), .B2(n162), .ZN(n17) );
  AOI22_X1 U18 ( .A1(a[3]), .A2(n159), .B1(b[3]), .B2(n156), .ZN(n18) );
  AOI22_X1 U19 ( .A1(a[0]), .A2(n157), .B1(b[0]), .B2(n154), .ZN(n68) );
  AOI22_X1 U20 ( .A1(a[1]), .A2(n157), .B1(b[1]), .B2(n154), .ZN(n46) );
  AOI22_X1 U21 ( .A1(a[2]), .A2(n158), .B1(b[2]), .B2(n155), .ZN(n24) );
  NAND2_X1 U22 ( .A1(n24), .A2(n25), .ZN(y[2]) );
  AOI22_X1 U23 ( .A1(c[2]), .A2(n164), .B1(d[2]), .B2(n161), .ZN(n25) );
  NAND2_X1 U24 ( .A1(n46), .A2(n47), .ZN(y[1]) );
  AOI22_X1 U25 ( .A1(c[1]), .A2(n163), .B1(d[1]), .B2(n160), .ZN(n47) );
  NAND2_X1 U26 ( .A1(n18), .A2(n19), .ZN(y[3]) );
  AOI22_X1 U27 ( .A1(c[3]), .A2(n165), .B1(d[3]), .B2(n162), .ZN(n19) );
  NAND2_X1 U28 ( .A1(n14), .A2(n15), .ZN(y[5]) );
  AOI22_X1 U29 ( .A1(a[5]), .A2(n159), .B1(b[5]), .B2(n156), .ZN(n14) );
  NAND2_X1 U30 ( .A1(n12), .A2(n13), .ZN(y[6]) );
  AOI22_X1 U31 ( .A1(a[6]), .A2(n159), .B1(b[6]), .B2(n156), .ZN(n12) );
  NAND2_X1 U32 ( .A1(n44), .A2(n45), .ZN(y[20]) );
  AOI22_X1 U33 ( .A1(a[20]), .A2(n158), .B1(b[20]), .B2(n155), .ZN(n44) );
  NAND2_X1 U34 ( .A1(n42), .A2(n43), .ZN(y[21]) );
  AOI22_X1 U35 ( .A1(a[21]), .A2(n158), .B1(b[21]), .B2(n155), .ZN(n42) );
  NAND2_X1 U36 ( .A1(n40), .A2(n41), .ZN(y[22]) );
  AOI22_X1 U37 ( .A1(a[22]), .A2(n158), .B1(b[22]), .B2(n155), .ZN(n40) );
  NAND2_X1 U38 ( .A1(n38), .A2(n39), .ZN(y[23]) );
  AOI22_X1 U39 ( .A1(a[23]), .A2(n158), .B1(b[23]), .B2(n155), .ZN(n38) );
  NAND2_X1 U40 ( .A1(n36), .A2(n37), .ZN(y[24]) );
  AOI22_X1 U41 ( .A1(a[24]), .A2(n158), .B1(b[24]), .B2(n155), .ZN(n36) );
  NAND2_X1 U42 ( .A1(n34), .A2(n35), .ZN(y[25]) );
  AOI22_X1 U43 ( .A1(a[25]), .A2(n158), .B1(b[25]), .B2(n155), .ZN(n34) );
  NAND2_X1 U44 ( .A1(n32), .A2(n33), .ZN(y[26]) );
  AOI22_X1 U45 ( .A1(a[26]), .A2(n158), .B1(b[26]), .B2(n155), .ZN(n32) );
  NAND2_X1 U46 ( .A1(n30), .A2(n31), .ZN(y[27]) );
  AOI22_X1 U47 ( .A1(a[27]), .A2(n158), .B1(b[27]), .B2(n155), .ZN(n30) );
  NAND2_X1 U48 ( .A1(n28), .A2(n29), .ZN(y[28]) );
  AOI22_X1 U49 ( .A1(a[28]), .A2(n158), .B1(b[28]), .B2(n155), .ZN(n28) );
  NAND2_X1 U50 ( .A1(n26), .A2(n27), .ZN(y[29]) );
  AOI22_X1 U51 ( .A1(a[29]), .A2(n158), .B1(b[29]), .B2(n155), .ZN(n26) );
  NAND2_X1 U52 ( .A1(n22), .A2(n23), .ZN(y[30]) );
  AOI22_X1 U53 ( .A1(a[30]), .A2(n158), .B1(b[30]), .B2(n155), .ZN(n22) );
  NAND2_X1 U54 ( .A1(n20), .A2(n21), .ZN(y[31]) );
  AOI22_X1 U55 ( .A1(a[31]), .A2(n159), .B1(b[31]), .B2(n156), .ZN(n20) );
  NAND2_X1 U56 ( .A1(n10), .A2(n11), .ZN(y[7]) );
  AOI22_X1 U57 ( .A1(a[7]), .A2(n159), .B1(b[7]), .B2(n156), .ZN(n10) );
  NAND2_X1 U58 ( .A1(n8), .A2(n9), .ZN(y[8]) );
  AOI22_X1 U59 ( .A1(a[8]), .A2(n159), .B1(b[8]), .B2(n156), .ZN(n8) );
  NAND2_X1 U60 ( .A1(n2), .A2(n3), .ZN(y[9]) );
  AOI22_X1 U61 ( .A1(a[9]), .A2(n159), .B1(b[9]), .B2(n156), .ZN(n2) );
  NAND2_X1 U62 ( .A1(n66), .A2(n67), .ZN(y[10]) );
  AOI22_X1 U63 ( .A1(a[10]), .A2(n157), .B1(b[10]), .B2(n154), .ZN(n66) );
  NAND2_X1 U64 ( .A1(n64), .A2(n65), .ZN(y[11]) );
  AOI22_X1 U65 ( .A1(a[11]), .A2(n157), .B1(b[11]), .B2(n154), .ZN(n64) );
  NAND2_X1 U66 ( .A1(n62), .A2(n63), .ZN(y[12]) );
  AOI22_X1 U67 ( .A1(a[12]), .A2(n157), .B1(b[12]), .B2(n154), .ZN(n62) );
  NAND2_X1 U68 ( .A1(n60), .A2(n61), .ZN(y[13]) );
  AOI22_X1 U69 ( .A1(a[13]), .A2(n157), .B1(b[13]), .B2(n154), .ZN(n60) );
  NAND2_X1 U70 ( .A1(n58), .A2(n59), .ZN(y[14]) );
  AOI22_X1 U71 ( .A1(a[14]), .A2(n157), .B1(b[14]), .B2(n154), .ZN(n58) );
  NAND2_X1 U72 ( .A1(n56), .A2(n57), .ZN(y[15]) );
  AOI22_X1 U73 ( .A1(a[15]), .A2(n157), .B1(b[15]), .B2(n154), .ZN(n56) );
  NAND2_X1 U74 ( .A1(n54), .A2(n55), .ZN(y[16]) );
  AOI22_X1 U75 ( .A1(a[16]), .A2(n157), .B1(b[16]), .B2(n154), .ZN(n54) );
  NAND2_X1 U76 ( .A1(n52), .A2(n53), .ZN(y[17]) );
  AOI22_X1 U77 ( .A1(a[17]), .A2(n157), .B1(b[17]), .B2(n154), .ZN(n52) );
  NAND2_X1 U78 ( .A1(n50), .A2(n51), .ZN(y[18]) );
  AOI22_X1 U79 ( .A1(a[18]), .A2(n157), .B1(b[18]), .B2(n154), .ZN(n50) );
  NAND2_X1 U80 ( .A1(n48), .A2(n49), .ZN(y[19]) );
  AOI22_X1 U81 ( .A1(a[19]), .A2(n157), .B1(b[19]), .B2(n154), .ZN(n48) );
  NOR2_X1 U82 ( .A1(sel[0]), .A2(sel[1]), .ZN(n6) );
  NOR2_X1 U83 ( .A1(n166), .A2(sel[1]), .ZN(n7) );
  AND2_X1 U84 ( .A1(sel[1]), .A2(n166), .ZN(n4) );
  AND2_X1 U85 ( .A1(sel[0]), .A2(sel[1]), .ZN(n5) );
  INV_X1 U86 ( .A(sel[0]), .ZN(n166) );
  AOI22_X1 U87 ( .A1(c[5]), .A2(n165), .B1(d[5]), .B2(n162), .ZN(n15) );
  AOI22_X1 U88 ( .A1(c[6]), .A2(n165), .B1(d[6]), .B2(n162), .ZN(n13) );
  AOI22_X1 U89 ( .A1(c[7]), .A2(n165), .B1(d[7]), .B2(n162), .ZN(n11) );
  AOI22_X1 U90 ( .A1(c[8]), .A2(n165), .B1(d[8]), .B2(n162), .ZN(n9) );
  AOI22_X1 U91 ( .A1(c[9]), .A2(n165), .B1(d[9]), .B2(n162), .ZN(n3) );
  AOI22_X1 U92 ( .A1(c[10]), .A2(n163), .B1(d[10]), .B2(n160), .ZN(n67) );
  AOI22_X1 U93 ( .A1(c[11]), .A2(n163), .B1(d[11]), .B2(n160), .ZN(n65) );
  AOI22_X1 U94 ( .A1(c[12]), .A2(n163), .B1(d[12]), .B2(n160), .ZN(n63) );
  AOI22_X1 U95 ( .A1(c[13]), .A2(n163), .B1(d[13]), .B2(n160), .ZN(n61) );
  AOI22_X1 U96 ( .A1(c[14]), .A2(n163), .B1(d[14]), .B2(n160), .ZN(n59) );
  AOI22_X1 U97 ( .A1(c[15]), .A2(n163), .B1(d[15]), .B2(n160), .ZN(n57) );
  AOI22_X1 U98 ( .A1(c[16]), .A2(n163), .B1(d[16]), .B2(n160), .ZN(n55) );
  AOI22_X1 U99 ( .A1(c[17]), .A2(n163), .B1(d[17]), .B2(n160), .ZN(n53) );
  AOI22_X1 U100 ( .A1(c[18]), .A2(n163), .B1(d[18]), .B2(n160), .ZN(n51) );
  AOI22_X1 U101 ( .A1(c[19]), .A2(n163), .B1(d[19]), .B2(n160), .ZN(n49) );
  AOI22_X1 U102 ( .A1(c[20]), .A2(n164), .B1(d[20]), .B2(n161), .ZN(n45) );
  AOI22_X1 U103 ( .A1(c[21]), .A2(n164), .B1(d[21]), .B2(n161), .ZN(n43) );
  AOI22_X1 U104 ( .A1(c[22]), .A2(n164), .B1(d[22]), .B2(n161), .ZN(n41) );
  AOI22_X1 U105 ( .A1(c[23]), .A2(n164), .B1(d[23]), .B2(n161), .ZN(n39) );
  AOI22_X1 U106 ( .A1(c[24]), .A2(n164), .B1(d[24]), .B2(n161), .ZN(n37) );
  AOI22_X1 U107 ( .A1(c[25]), .A2(n164), .B1(d[25]), .B2(n161), .ZN(n35) );
  AOI22_X1 U108 ( .A1(c[26]), .A2(n164), .B1(d[26]), .B2(n161), .ZN(n33) );
  AOI22_X1 U109 ( .A1(c[27]), .A2(n164), .B1(d[27]), .B2(n161), .ZN(n31) );
  AOI22_X1 U110 ( .A1(c[28]), .A2(n164), .B1(d[28]), .B2(n161), .ZN(n29) );
  AOI22_X1 U111 ( .A1(c[29]), .A2(n164), .B1(d[29]), .B2(n161), .ZN(n27) );
  AOI22_X1 U112 ( .A1(c[30]), .A2(n164), .B1(d[30]), .B2(n161), .ZN(n23) );
  AOI22_X1 U113 ( .A1(c[31]), .A2(n165), .B1(d[31]), .B2(n162), .ZN(n21) );
endmodule


module Mux21_5 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148;

  BUF_X1 U1 ( .A(n148), .Z(n140) );
  BUF_X1 U2 ( .A(n145), .Z(n147) );
  BUF_X1 U3 ( .A(n143), .Z(n146) );
  BUF_X1 U4 ( .A(n148), .Z(n145) );
  BUF_X1 U5 ( .A(n148), .Z(n144) );
  BUF_X1 U6 ( .A(n148), .Z(n141) );
  BUF_X1 U7 ( .A(n148), .Z(n143) );
  BUF_X1 U8 ( .A(n148), .Z(n142) );
  INV_X1 U9 ( .A(n139), .ZN(n148) );
  INV_X1 U10 ( .A(n38), .ZN(y[5]) );
  AOI22_X1 U11 ( .A1(a[5]), .A2(sel), .B1(b[5]), .B2(n141), .ZN(n38) );
  INV_X1 U12 ( .A(n37), .ZN(y[6]) );
  AOI22_X1 U13 ( .A1(a[6]), .A2(n139), .B1(b[6]), .B2(n140), .ZN(n37) );
  INV_X1 U14 ( .A(n62), .ZN(y[12]) );
  AOI22_X1 U15 ( .A1(a[12]), .A2(sel), .B1(b[12]), .B2(n147), .ZN(n62) );
  INV_X1 U16 ( .A(n61), .ZN(y[13]) );
  AOI22_X1 U17 ( .A1(a[13]), .A2(n139), .B1(b[13]), .B2(n146), .ZN(n61) );
  INV_X1 U18 ( .A(n60), .ZN(y[14]) );
  AOI22_X1 U19 ( .A1(a[14]), .A2(sel), .B1(b[14]), .B2(n146), .ZN(n60) );
  INV_X1 U20 ( .A(n34), .ZN(y[9]) );
  AOI22_X1 U21 ( .A1(n139), .A2(a[9]), .B1(b[9]), .B2(n140), .ZN(n34) );
  INV_X1 U22 ( .A(n35), .ZN(y[8]) );
  AOI22_X1 U23 ( .A1(a[8]), .A2(sel), .B1(b[8]), .B2(n140), .ZN(n35) );
  INV_X1 U24 ( .A(n39), .ZN(y[4]) );
  AOI22_X1 U25 ( .A1(a[4]), .A2(n139), .B1(b[4]), .B2(n141), .ZN(n39) );
  INV_X1 U26 ( .A(n40), .ZN(y[3]) );
  AOI22_X1 U27 ( .A1(a[3]), .A2(sel), .B1(b[3]), .B2(n141), .ZN(n40) );
  INV_X1 U28 ( .A(n43), .ZN(y[2]) );
  AOI22_X1 U29 ( .A1(a[2]), .A2(sel), .B1(b[2]), .B2(n142), .ZN(n43) );
  INV_X1 U30 ( .A(n36), .ZN(y[7]) );
  AOI22_X1 U31 ( .A1(a[7]), .A2(n139), .B1(b[7]), .B2(n140), .ZN(n36) );
  INV_X1 U32 ( .A(n64), .ZN(y[10]) );
  AOI22_X1 U33 ( .A1(a[10]), .A2(n139), .B1(b[10]), .B2(n147), .ZN(n64) );
  INV_X1 U34 ( .A(n63), .ZN(y[11]) );
  AOI22_X1 U35 ( .A1(a[11]), .A2(sel), .B1(b[11]), .B2(n147), .ZN(n63) );
  INV_X1 U36 ( .A(n65), .ZN(y[0]) );
  AOI22_X1 U37 ( .A1(a[0]), .A2(n139), .B1(b[0]), .B2(n147), .ZN(n65) );
  INV_X1 U38 ( .A(n51), .ZN(y[22]) );
  INV_X1 U39 ( .A(n48), .ZN(y[25]) );
  INV_X1 U40 ( .A(n47), .ZN(y[26]) );
  INV_X1 U41 ( .A(n46), .ZN(y[27]) );
  INV_X1 U42 ( .A(n45), .ZN(y[28]) );
  INV_X1 U43 ( .A(n44), .ZN(y[29]) );
  INV_X1 U44 ( .A(n42), .ZN(y[30]) );
  INV_X1 U45 ( .A(n41), .ZN(y[31]) );
  INV_X1 U46 ( .A(n59), .ZN(y[15]) );
  AOI22_X1 U47 ( .A1(a[15]), .A2(sel), .B1(b[15]), .B2(n146), .ZN(n59) );
  INV_X1 U48 ( .A(n58), .ZN(y[16]) );
  AOI22_X1 U49 ( .A1(a[16]), .A2(n139), .B1(b[16]), .B2(n146), .ZN(n58) );
  INV_X1 U50 ( .A(n57), .ZN(y[17]) );
  AOI22_X1 U51 ( .A1(a[17]), .A2(sel), .B1(b[17]), .B2(n145), .ZN(n57) );
  INV_X1 U52 ( .A(n56), .ZN(y[18]) );
  AOI22_X1 U53 ( .A1(a[18]), .A2(n139), .B1(b[18]), .B2(n145), .ZN(n56) );
  INV_X1 U54 ( .A(n55), .ZN(y[19]) );
  AOI22_X1 U55 ( .A1(a[19]), .A2(sel), .B1(b[19]), .B2(n145), .ZN(n55) );
  INV_X1 U56 ( .A(n53), .ZN(y[20]) );
  AOI22_X1 U57 ( .A1(a[20]), .A2(n139), .B1(b[20]), .B2(n144), .ZN(n53) );
  INV_X1 U58 ( .A(n52), .ZN(y[21]) );
  AOI22_X1 U59 ( .A1(a[21]), .A2(sel), .B1(b[21]), .B2(n144), .ZN(n52) );
  INV_X1 U60 ( .A(n50), .ZN(y[23]) );
  AOI22_X1 U61 ( .A1(a[23]), .A2(n139), .B1(b[23]), .B2(n144), .ZN(n50) );
  INV_X1 U62 ( .A(n49), .ZN(y[24]) );
  AOI22_X1 U63 ( .A1(a[24]), .A2(sel), .B1(b[24]), .B2(n143), .ZN(n49) );
  INV_X1 U64 ( .A(n54), .ZN(y[1]) );
  AOI22_X1 U65 ( .A1(a[1]), .A2(n139), .B1(b[1]), .B2(n145), .ZN(n54) );
  BUF_X1 U66 ( .A(sel), .Z(n139) );
  AOI22_X1 U67 ( .A1(a[22]), .A2(n139), .B1(b[22]), .B2(n144), .ZN(n51) );
  AOI22_X1 U68 ( .A1(a[31]), .A2(sel), .B1(b[31]), .B2(n141), .ZN(n41) );
  AOI22_X1 U69 ( .A1(a[30]), .A2(n139), .B1(b[30]), .B2(n142), .ZN(n42) );
  AOI22_X1 U70 ( .A1(a[29]), .A2(sel), .B1(b[29]), .B2(n142), .ZN(n44) );
  AOI22_X1 U71 ( .A1(a[28]), .A2(n139), .B1(b[28]), .B2(n142), .ZN(n45) );
  AOI22_X1 U72 ( .A1(a[27]), .A2(sel), .B1(b[27]), .B2(n143), .ZN(n46) );
  AOI22_X1 U73 ( .A1(a[26]), .A2(n139), .B1(b[26]), .B2(n143), .ZN(n47) );
  AOI22_X1 U74 ( .A1(a[25]), .A2(sel), .B1(b[25]), .B2(n143), .ZN(n48) );
endmodule


module BranchUnit ( a, sel, y );
  input [31:0] a;
  input sel;
  output y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;

  NOR4_X1 U2 ( .A1(a[5]), .A2(a[4]), .A3(a[3]), .A4(a[31]), .ZN(n10) );
  NOR4_X1 U3 ( .A1(a[1]), .A2(a[19]), .A3(a[18]), .A4(a[17]), .ZN(n6) );
  NOR4_X1 U4 ( .A1(a[12]), .A2(a[11]), .A3(a[10]), .A4(a[0]), .ZN(n4) );
  NOR4_X1 U5 ( .A1(a[16]), .A2(a[15]), .A3(a[14]), .A4(a[13]), .ZN(n5) );
  NOR4_X1 U6 ( .A1(a[30]), .A2(a[2]), .A3(a[29]), .A4(a[28]), .ZN(n9) );
  NOR4_X1 U7 ( .A1(a[27]), .A2(a[26]), .A3(a[25]), .A4(a[24]), .ZN(n8) );
  NOR2_X1 U8 ( .A1(n2), .A2(n3), .ZN(n1) );
  NAND4_X1 U9 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n2) );
  NOR4_X1 U10 ( .A1(a[9]), .A2(a[8]), .A3(a[7]), .A4(a[6]), .ZN(n11) );
  NAND4_X1 U11 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(n3) );
  NOR4_X1 U12 ( .A1(a[23]), .A2(a[22]), .A3(a[21]), .A4(a[20]), .ZN(n7) );
  XNOR2_X1 U13 ( .A(sel), .B(n1), .ZN(y) );
endmodule


module reg_11 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n177) );
  BUF_X1 U4 ( .A(n35), .Z(n176) );
  BUF_X1 U5 ( .A(n35), .Z(n178) );
  BUF_X1 U6 ( .A(n34), .Z(n179) );
  BUF_X1 U7 ( .A(n34), .Z(n180) );
  BUF_X1 U8 ( .A(n34), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n35) );
  OAI22_X1 U10 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U11 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U12 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U13 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U14 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U15 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U16 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U17 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U18 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U19 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U20 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U21 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U22 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U23 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U24 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U25 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U26 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U27 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U28 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n205) );
  OAI22_X1 U30 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U31 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U32 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U33 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U34 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U35 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U36 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U37 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U38 ( .A1(n179), .A2(n58), .B1(n176), .B2(n185), .ZN(n77) );
  INV_X1 U39 ( .A(i[22]), .ZN(n185) );
  OAI22_X1 U40 ( .A1(n179), .A2(n61), .B1(n176), .B2(n193), .ZN(n74) );
  INV_X1 U41 ( .A(i[25]), .ZN(n193) );
  OAI22_X1 U42 ( .A1(n179), .A2(n62), .B1(n176), .B2(n194), .ZN(n73) );
  INV_X1 U43 ( .A(i[26]), .ZN(n194) );
  OAI22_X1 U44 ( .A1(n179), .A2(n63), .B1(n176), .B2(n195), .ZN(n72) );
  INV_X1 U45 ( .A(i[27]), .ZN(n195) );
  OAI22_X1 U46 ( .A1(n179), .A2(n64), .B1(n176), .B2(n196), .ZN(n71) );
  INV_X1 U47 ( .A(i[28]), .ZN(n196) );
  OAI22_X1 U48 ( .A1(n179), .A2(n65), .B1(n176), .B2(n197), .ZN(n70) );
  INV_X1 U49 ( .A(i[29]), .ZN(n197) );
  OAI22_X1 U50 ( .A1(n179), .A2(n66), .B1(n176), .B2(n198), .ZN(n69) );
  INV_X1 U51 ( .A(i[30]), .ZN(n198) );
  OAI22_X1 U52 ( .A1(n179), .A2(n67), .B1(n176), .B2(n199), .ZN(n68) );
  INV_X1 U53 ( .A(i[31]), .ZN(n199) );
  OAI22_X1 U54 ( .A1(n180), .A2(n51), .B1(n177), .B2(n192), .ZN(n84) );
  INV_X1 U55 ( .A(i[15]), .ZN(n192) );
  OAI22_X1 U56 ( .A1(n180), .A2(n52), .B1(n177), .B2(n191), .ZN(n83) );
  INV_X1 U57 ( .A(i[16]), .ZN(n191) );
  OAI22_X1 U58 ( .A1(n180), .A2(n53), .B1(n177), .B2(n190), .ZN(n82) );
  INV_X1 U59 ( .A(i[17]), .ZN(n190) );
  OAI22_X1 U60 ( .A1(n180), .A2(n54), .B1(n177), .B2(n189), .ZN(n81) );
  INV_X1 U61 ( .A(i[18]), .ZN(n189) );
  OAI22_X1 U62 ( .A1(n180), .A2(n55), .B1(n177), .B2(n188), .ZN(n80) );
  INV_X1 U63 ( .A(i[19]), .ZN(n188) );
  OAI22_X1 U64 ( .A1(n179), .A2(n56), .B1(n176), .B2(n187), .ZN(n79) );
  INV_X1 U65 ( .A(i[20]), .ZN(n187) );
  OAI22_X1 U66 ( .A1(n179), .A2(n57), .B1(n176), .B2(n186), .ZN(n78) );
  INV_X1 U67 ( .A(i[21]), .ZN(n186) );
  OAI22_X1 U68 ( .A1(n179), .A2(n59), .B1(n176), .B2(n184), .ZN(n76) );
  INV_X1 U69 ( .A(i[23]), .ZN(n184) );
  OAI22_X1 U70 ( .A1(n179), .A2(n60), .B1(n176), .B2(n183), .ZN(n75) );
  INV_X1 U71 ( .A(i[24]), .ZN(n183) );
  OAI22_X1 U72 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U73 ( .A(i[1]), .ZN(n213) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n34) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module reg_10 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n177) );
  BUF_X1 U4 ( .A(n35), .Z(n176) );
  BUF_X1 U5 ( .A(n35), .Z(n178) );
  BUF_X1 U6 ( .A(n34), .Z(n179) );
  BUF_X1 U7 ( .A(n34), .Z(n180) );
  BUF_X1 U8 ( .A(n34), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n35) );
  OAI22_X1 U10 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U11 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U12 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U13 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U14 ( .A1(n180), .A2(n52), .B1(n177), .B2(n198), .ZN(n83) );
  INV_X1 U15 ( .A(i[16]), .ZN(n198) );
  OAI22_X1 U16 ( .A1(n179), .A2(n56), .B1(n176), .B2(n194), .ZN(n79) );
  INV_X1 U17 ( .A(i[20]), .ZN(n194) );
  OAI22_X1 U18 ( .A1(n179), .A2(n63), .B1(n176), .B2(n187), .ZN(n72) );
  INV_X1 U19 ( .A(i[27]), .ZN(n187) );
  OAI22_X1 U20 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U21 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U22 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U23 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U24 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U25 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U26 ( .A1(n180), .A2(n53), .B1(n177), .B2(n197), .ZN(n82) );
  INV_X1 U27 ( .A(i[17]), .ZN(n197) );
  OAI22_X1 U28 ( .A1(n179), .A2(n60), .B1(n176), .B2(n190), .ZN(n75) );
  INV_X1 U29 ( .A(i[24]), .ZN(n190) );
  OAI22_X1 U30 ( .A1(n179), .A2(n64), .B1(n176), .B2(n186), .ZN(n71) );
  INV_X1 U31 ( .A(i[28]), .ZN(n186) );
  OAI22_X1 U32 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U33 ( .A(i[31]), .ZN(n183) );
  OAI22_X1 U34 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U35 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U36 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U37 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U38 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U40 ( .A1(n180), .A2(n54), .B1(n177), .B2(n196), .ZN(n81) );
  INV_X1 U41 ( .A(i[18]), .ZN(n196) );
  OAI22_X1 U42 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U43 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U44 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U45 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U46 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U47 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U48 ( .A1(n179), .A2(n57), .B1(n176), .B2(n193), .ZN(n78) );
  INV_X1 U49 ( .A(i[21]), .ZN(n193) );
  OAI22_X1 U50 ( .A1(n179), .A2(n61), .B1(n176), .B2(n189), .ZN(n74) );
  INV_X1 U51 ( .A(i[25]), .ZN(n189) );
  OAI22_X1 U52 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U53 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U54 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U55 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U56 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U57 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U58 ( .A1(n180), .A2(n51), .B1(n177), .B2(n199), .ZN(n84) );
  INV_X1 U59 ( .A(i[15]), .ZN(n199) );
  OAI22_X1 U60 ( .A1(n180), .A2(n55), .B1(n177), .B2(n195), .ZN(n80) );
  INV_X1 U61 ( .A(i[19]), .ZN(n195) );
  OAI22_X1 U62 ( .A1(n179), .A2(n62), .B1(n176), .B2(n188), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n188) );
  OAI22_X1 U64 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U65 ( .A(i[1]), .ZN(n213) );
  OAI22_X1 U66 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U67 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U68 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U69 ( .A(i[9]), .ZN(n205) );
  OAI22_X1 U70 ( .A1(n179), .A2(n59), .B1(n176), .B2(n191), .ZN(n76) );
  INV_X1 U71 ( .A(i[23]), .ZN(n191) );
  OAI22_X1 U72 ( .A1(n179), .A2(n58), .B1(n176), .B2(n192), .ZN(n77) );
  INV_X1 U73 ( .A(i[22]), .ZN(n192) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n34) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module reg_9 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n34, n35, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n35), .Z(n177) );
  BUF_X1 U4 ( .A(n35), .Z(n176) );
  BUF_X1 U5 ( .A(n35), .Z(n178) );
  BUF_X1 U6 ( .A(n34), .Z(n179) );
  BUF_X1 U7 ( .A(n34), .Z(n180) );
  BUF_X1 U8 ( .A(n34), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n35) );
  OAI22_X1 U10 ( .A1(n179), .A2(n60), .B1(n176), .B2(n190), .ZN(n75) );
  INV_X1 U11 ( .A(i[24]), .ZN(n190) );
  OAI22_X1 U12 ( .A1(n179), .A2(n61), .B1(n176), .B2(n189), .ZN(n74) );
  INV_X1 U13 ( .A(i[25]), .ZN(n189) );
  OAI22_X1 U14 ( .A1(n179), .A2(n62), .B1(n176), .B2(n188), .ZN(n73) );
  INV_X1 U15 ( .A(i[26]), .ZN(n188) );
  OAI22_X1 U16 ( .A1(n179), .A2(n63), .B1(n176), .B2(n187), .ZN(n72) );
  INV_X1 U17 ( .A(i[27]), .ZN(n187) );
  OAI22_X1 U18 ( .A1(n179), .A2(n64), .B1(n176), .B2(n186), .ZN(n71) );
  INV_X1 U19 ( .A(i[28]), .ZN(n186) );
  OAI22_X1 U20 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U21 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U22 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U23 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U24 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U25 ( .A(i[31]), .ZN(n183) );
  OAI22_X1 U26 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U27 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U28 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U29 ( .A(i[1]), .ZN(n213) );
  OAI22_X1 U30 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U31 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U32 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U33 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U34 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U35 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U36 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U37 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U38 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U39 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U40 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U41 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U42 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U43 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U44 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U45 ( .A(i[9]), .ZN(n205) );
  OAI22_X1 U46 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U47 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U48 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U49 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U50 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U51 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U52 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U53 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U54 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U55 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U56 ( .A1(n180), .A2(n51), .B1(n177), .B2(n199), .ZN(n84) );
  INV_X1 U57 ( .A(i[15]), .ZN(n199) );
  OAI22_X1 U58 ( .A1(n180), .A2(n52), .B1(n177), .B2(n198), .ZN(n83) );
  INV_X1 U59 ( .A(i[16]), .ZN(n198) );
  OAI22_X1 U60 ( .A1(n180), .A2(n53), .B1(n177), .B2(n197), .ZN(n82) );
  INV_X1 U61 ( .A(i[17]), .ZN(n197) );
  OAI22_X1 U62 ( .A1(n180), .A2(n54), .B1(n177), .B2(n196), .ZN(n81) );
  INV_X1 U63 ( .A(i[18]), .ZN(n196) );
  OAI22_X1 U64 ( .A1(n180), .A2(n55), .B1(n177), .B2(n195), .ZN(n80) );
  INV_X1 U65 ( .A(i[19]), .ZN(n195) );
  OAI22_X1 U66 ( .A1(n179), .A2(n56), .B1(n176), .B2(n194), .ZN(n79) );
  INV_X1 U67 ( .A(i[20]), .ZN(n194) );
  OAI22_X1 U68 ( .A1(n179), .A2(n57), .B1(n176), .B2(n193), .ZN(n78) );
  INV_X1 U69 ( .A(i[21]), .ZN(n193) );
  OAI22_X1 U70 ( .A1(n179), .A2(n58), .B1(n176), .B2(n192), .ZN(n77) );
  INV_X1 U71 ( .A(i[22]), .ZN(n192) );
  OAI22_X1 U72 ( .A1(n179), .A2(n59), .B1(n176), .B2(n191), .ZN(n76) );
  INV_X1 U73 ( .A(i[23]), .ZN(n191) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n34) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module reg_8 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n215), .Z(n177) );
  BUF_X1 U4 ( .A(n215), .Z(n176) );
  BUF_X1 U5 ( .A(n215), .Z(n178) );
  BUF_X1 U6 ( .A(n216), .Z(n179) );
  BUF_X1 U7 ( .A(n216), .Z(n180) );
  BUF_X1 U8 ( .A(n216), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n215) );
  OAI22_X1 U10 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U11 ( .A(i[1]), .ZN(n213) );
  OAI22_X1 U12 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U13 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U14 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U15 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U16 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U17 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U18 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U19 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U20 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U21 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U22 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U23 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U24 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U25 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U26 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U27 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U28 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U29 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U30 ( .A1(n180), .A2(n51), .B1(n177), .B2(n199), .ZN(n84) );
  INV_X1 U31 ( .A(i[15]), .ZN(n199) );
  OAI22_X1 U32 ( .A1(n180), .A2(n52), .B1(n177), .B2(n198), .ZN(n83) );
  INV_X1 U33 ( .A(i[16]), .ZN(n198) );
  OAI22_X1 U34 ( .A1(n180), .A2(n53), .B1(n177), .B2(n197), .ZN(n82) );
  INV_X1 U35 ( .A(i[17]), .ZN(n197) );
  OAI22_X1 U36 ( .A1(n180), .A2(n54), .B1(n177), .B2(n196), .ZN(n81) );
  INV_X1 U37 ( .A(i[18]), .ZN(n196) );
  OAI22_X1 U38 ( .A1(n180), .A2(n55), .B1(n177), .B2(n195), .ZN(n80) );
  INV_X1 U39 ( .A(i[19]), .ZN(n195) );
  OAI22_X1 U40 ( .A1(n179), .A2(n56), .B1(n176), .B2(n194), .ZN(n79) );
  INV_X1 U41 ( .A(i[20]), .ZN(n194) );
  OAI22_X1 U42 ( .A1(n179), .A2(n57), .B1(n176), .B2(n193), .ZN(n78) );
  INV_X1 U43 ( .A(i[21]), .ZN(n193) );
  OAI22_X1 U44 ( .A1(n179), .A2(n58), .B1(n176), .B2(n192), .ZN(n77) );
  INV_X1 U45 ( .A(i[22]), .ZN(n192) );
  OAI22_X1 U46 ( .A1(n179), .A2(n59), .B1(n176), .B2(n191), .ZN(n76) );
  INV_X1 U47 ( .A(i[23]), .ZN(n191) );
  OAI22_X1 U48 ( .A1(n179), .A2(n60), .B1(n176), .B2(n190), .ZN(n75) );
  INV_X1 U49 ( .A(i[24]), .ZN(n190) );
  OAI22_X1 U50 ( .A1(n179), .A2(n61), .B1(n176), .B2(n189), .ZN(n74) );
  INV_X1 U51 ( .A(i[25]), .ZN(n189) );
  OAI22_X1 U52 ( .A1(n179), .A2(n62), .B1(n176), .B2(n188), .ZN(n73) );
  INV_X1 U53 ( .A(i[26]), .ZN(n188) );
  OAI22_X1 U54 ( .A1(n179), .A2(n63), .B1(n176), .B2(n187), .ZN(n72) );
  INV_X1 U55 ( .A(i[27]), .ZN(n187) );
  OAI22_X1 U56 ( .A1(n179), .A2(n64), .B1(n176), .B2(n186), .ZN(n71) );
  INV_X1 U57 ( .A(i[28]), .ZN(n186) );
  OAI22_X1 U58 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U59 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U60 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U61 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U62 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U63 ( .A(i[31]), .ZN(n183) );
  OAI22_X1 U64 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U65 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U66 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U67 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U68 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U69 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U70 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U71 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U72 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U73 ( .A(i[9]), .ZN(n205) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n216) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module reg_7 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n215), .Z(n177) );
  BUF_X1 U4 ( .A(n215), .Z(n176) );
  BUF_X1 U5 ( .A(n215), .Z(n178) );
  BUF_X1 U6 ( .A(n216), .Z(n179) );
  BUF_X1 U7 ( .A(n216), .Z(n180) );
  BUF_X1 U8 ( .A(n216), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n215) );
  OAI22_X1 U10 ( .A1(n181), .A2(n36), .B1(n178), .B2(n187), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n187) );
  OAI22_X1 U12 ( .A1(n181), .A2(n40), .B1(n178), .B2(n183), .ZN(n95) );
  INV_X1 U13 ( .A(i[4]), .ZN(n183) );
  OAI22_X1 U14 ( .A1(n181), .A2(n38), .B1(n178), .B2(n185), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n185) );
  OAI22_X1 U16 ( .A1(n181), .A2(n37), .B1(n178), .B2(n186), .ZN(n98) );
  INV_X1 U17 ( .A(i[1]), .ZN(n186) );
  OAI22_X1 U18 ( .A1(n181), .A2(n39), .B1(n178), .B2(n184), .ZN(n96) );
  INV_X1 U19 ( .A(i[3]), .ZN(n184) );
  OAI22_X1 U20 ( .A1(n181), .A2(n41), .B1(n178), .B2(n188), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n188) );
  OAI22_X1 U22 ( .A1(n181), .A2(n42), .B1(n178), .B2(n189), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n189) );
  OAI22_X1 U24 ( .A1(n179), .A2(n56), .B1(n176), .B2(n203), .ZN(n79) );
  INV_X1 U25 ( .A(i[20]), .ZN(n203) );
  OAI22_X1 U26 ( .A1(n179), .A2(n57), .B1(n176), .B2(n204), .ZN(n78) );
  INV_X1 U27 ( .A(i[21]), .ZN(n204) );
  OAI22_X1 U28 ( .A1(n179), .A2(n58), .B1(n176), .B2(n205), .ZN(n77) );
  INV_X1 U29 ( .A(i[22]), .ZN(n205) );
  OAI22_X1 U30 ( .A1(n179), .A2(n59), .B1(n176), .B2(n206), .ZN(n76) );
  INV_X1 U31 ( .A(i[23]), .ZN(n206) );
  OAI22_X1 U32 ( .A1(n179), .A2(n60), .B1(n176), .B2(n207), .ZN(n75) );
  INV_X1 U33 ( .A(i[24]), .ZN(n207) );
  OAI22_X1 U34 ( .A1(n179), .A2(n61), .B1(n176), .B2(n208), .ZN(n74) );
  INV_X1 U35 ( .A(i[25]), .ZN(n208) );
  OAI22_X1 U36 ( .A1(n179), .A2(n62), .B1(n176), .B2(n209), .ZN(n73) );
  INV_X1 U37 ( .A(i[26]), .ZN(n209) );
  OAI22_X1 U38 ( .A1(n179), .A2(n63), .B1(n176), .B2(n210), .ZN(n72) );
  INV_X1 U39 ( .A(i[27]), .ZN(n210) );
  OAI22_X1 U40 ( .A1(n179), .A2(n64), .B1(n176), .B2(n211), .ZN(n71) );
  INV_X1 U41 ( .A(i[28]), .ZN(n211) );
  OAI22_X1 U42 ( .A1(n179), .A2(n65), .B1(n176), .B2(n212), .ZN(n70) );
  INV_X1 U43 ( .A(i[29]), .ZN(n212) );
  OAI22_X1 U44 ( .A1(n179), .A2(n66), .B1(n176), .B2(n213), .ZN(n69) );
  INV_X1 U45 ( .A(i[30]), .ZN(n213) );
  OAI22_X1 U46 ( .A1(n179), .A2(n67), .B1(n176), .B2(n214), .ZN(n68) );
  INV_X1 U47 ( .A(i[31]), .ZN(n214) );
  OAI22_X1 U48 ( .A1(n180), .A2(n43), .B1(n178), .B2(n190), .ZN(n92) );
  INV_X1 U49 ( .A(i[7]), .ZN(n190) );
  OAI22_X1 U50 ( .A1(n180), .A2(n44), .B1(n177), .B2(n191), .ZN(n91) );
  INV_X1 U51 ( .A(i[8]), .ZN(n191) );
  OAI22_X1 U52 ( .A1(n180), .A2(n45), .B1(n177), .B2(n192), .ZN(n90) );
  INV_X1 U53 ( .A(i[9]), .ZN(n192) );
  OAI22_X1 U54 ( .A1(n180), .A2(n46), .B1(n177), .B2(n193), .ZN(n89) );
  INV_X1 U55 ( .A(i[10]), .ZN(n193) );
  OAI22_X1 U56 ( .A1(n180), .A2(n47), .B1(n177), .B2(n194), .ZN(n88) );
  INV_X1 U57 ( .A(i[11]), .ZN(n194) );
  OAI22_X1 U58 ( .A1(n180), .A2(n48), .B1(n177), .B2(n195), .ZN(n87) );
  INV_X1 U59 ( .A(i[12]), .ZN(n195) );
  OAI22_X1 U60 ( .A1(n180), .A2(n49), .B1(n177), .B2(n196), .ZN(n86) );
  INV_X1 U61 ( .A(i[13]), .ZN(n196) );
  OAI22_X1 U62 ( .A1(n180), .A2(n50), .B1(n177), .B2(n197), .ZN(n85) );
  INV_X1 U63 ( .A(i[14]), .ZN(n197) );
  OAI22_X1 U64 ( .A1(n180), .A2(n51), .B1(n177), .B2(n198), .ZN(n84) );
  INV_X1 U65 ( .A(i[15]), .ZN(n198) );
  OAI22_X1 U66 ( .A1(n180), .A2(n52), .B1(n177), .B2(n199), .ZN(n83) );
  INV_X1 U67 ( .A(i[16]), .ZN(n199) );
  OAI22_X1 U68 ( .A1(n180), .A2(n53), .B1(n177), .B2(n200), .ZN(n82) );
  INV_X1 U69 ( .A(i[17]), .ZN(n200) );
  OAI22_X1 U70 ( .A1(n180), .A2(n54), .B1(n177), .B2(n201), .ZN(n81) );
  INV_X1 U71 ( .A(i[18]), .ZN(n201) );
  OAI22_X1 U72 ( .A1(n180), .A2(n55), .B1(n177), .B2(n202), .ZN(n80) );
  INV_X1 U73 ( .A(i[19]), .ZN(n202) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n216) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module register_file ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, ADD_RD1, 
        ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700,
         N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711,
         N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N1020,
         N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030,
         N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040,
         N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050,
         N1051, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3448,
         n3450, n3452, n3453, n3456, n3458, n3459, n3460, n3461, n3462, n3464,
         n3466, n3468, n3469, n3472, n3474, n3475, n3476, n3477, n3478, n3480,
         n3482, n3484, n3485, n3488, n3490, n3491, n3492, n3493, n3494, n3496,
         n3498, n3500, n3501, n3504, n3506, n3507, n3508, n3509, n3510, n3512,
         n3514, n3516, n3517, n3520, n3522, n3523, n3524, n3525, n3526, n3528,
         n3530, n3532, n3533, n3536, n3538, n3539, n3540, n3541, n3542, n3544,
         n3546, n3548, n3549, n3552, n3554, n3555, n3556, n3557, n3558, n3560,
         n3562, n3564, n3565, n3568, n3570, n3571, n3572, n3573, n3574, n3576,
         n3578, n3580, n3581, n3584, n3586, n3587, n3588, n3589, n3590, n3592,
         n3594, n3596, n3597, n3600, n3602, n3603, n3604, n3605, n3606, n3608,
         n3610, n3612, n3613, n3616, n3618, n3619, n3620, n3621, n3622, n3624,
         n3626, n3628, n3629, n3632, n3634, n3635, n3636, n3637, n3638, n3640,
         n3642, n3644, n3645, n3648, n3650, n3651, n3652, n3653, n3654, n3656,
         n3658, n3660, n3661, n3664, n3666, n3667, n3668, n3669, n3670, n3672,
         n3674, n3676, n3677, n3680, n3682, n3683, n3684, n3685, n3686, n3688,
         n3690, n3692, n3693, n3696, n3698, n3699, n3700, n3701, n3702, n3704,
         n3706, n3708, n3709, n3712, n3714, n3715, n3716, n3717, n3718, n3720,
         n3722, n3724, n3725, n3728, n3730, n3731, n3732, n3733, n3734, n3736,
         n3738, n3740, n3741, n3744, n3746, n3747, n3748, n3749, n3750, n3752,
         n3754, n3756, n3757, n3760, n3762, n3763, n3764, n3765, n3766, n3768,
         n3770, n3772, n3773, n3776, n3778, n3779, n3780, n3781, n3782, n3784,
         n3786, n3788, n3789, n3792, n3794, n3795, n3796, n3797, n3798, n3800,
         n3802, n3804, n3805, n3808, n3810, n3811, n3812, n3813, n3814, n3816,
         n3818, n3820, n3821, n3824, n3826, n3827, n3828, n3829, n3830, n3832,
         n3834, n3836, n3837, n3840, n3842, n3843, n3844, n3845, n3846, n3848,
         n3850, n3852, n3853, n3856, n3858, n3859, n3860, n3861, n3862, n3864,
         n3866, n3868, n3869, n3872, n3874, n3875, n3876, n3877, n3878, n3880,
         n3882, n3884, n3885, n3888, n3890, n3891, n3892, n3893, n3894, n3896,
         n3898, n3900, n3901, n3904, n3906, n3907, n3908, n3909, n3910, n3912,
         n3914, n3916, n3917, n3920, n3922, n3923, n3924, n3925, n3926, n3928,
         n3930, n3932, n3933, n3936, n3938, n3939, n3940, n3941, n3942, n3944,
         n3946, n3948, n3949, n3952, n3954, n3955, n3956, n3957, n3958, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n815, n816, n817, n819, n821, n822, n824, n826,
         n827, n830, n842, n845, n847, n849, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665;
  assign OUT1[0] = N690;
  assign OUT1[1] = N691;
  assign OUT1[2] = N692;
  assign OUT1[3] = N693;
  assign OUT1[4] = N694;
  assign OUT1[5] = N695;
  assign OUT1[6] = N696;
  assign OUT1[7] = N697;
  assign OUT1[8] = N698;
  assign OUT1[9] = N699;
  assign OUT1[10] = N700;
  assign OUT1[11] = N701;
  assign OUT1[12] = N702;
  assign OUT1[13] = N703;
  assign OUT1[14] = N704;
  assign OUT1[15] = N705;
  assign OUT1[16] = N706;
  assign OUT1[17] = N707;
  assign OUT1[18] = N708;
  assign OUT1[19] = N709;
  assign OUT1[20] = N710;
  assign OUT1[21] = N711;
  assign OUT1[22] = N712;
  assign OUT1[23] = N713;
  assign OUT1[24] = N714;
  assign OUT1[25] = N715;
  assign OUT1[26] = N716;
  assign OUT1[27] = N717;
  assign OUT1[28] = N718;
  assign OUT1[29] = N719;
  assign OUT1[30] = N720;
  assign OUT1[31] = N721;
  assign OUT2[0] = N1020;
  assign OUT2[1] = N1021;
  assign OUT2[2] = N1022;
  assign OUT2[3] = N1023;
  assign OUT2[4] = N1024;
  assign OUT2[5] = N1025;
  assign OUT2[6] = N1026;
  assign OUT2[7] = N1027;
  assign OUT2[8] = N1028;
  assign OUT2[9] = N1029;
  assign OUT2[10] = N1030;
  assign OUT2[11] = N1031;
  assign OUT2[12] = N1032;
  assign OUT2[13] = N1033;
  assign OUT2[14] = N1034;
  assign OUT2[15] = N1035;
  assign OUT2[16] = N1036;
  assign OUT2[17] = N1037;
  assign OUT2[18] = N1038;
  assign OUT2[19] = N1039;
  assign OUT2[20] = N1040;
  assign OUT2[21] = N1041;
  assign OUT2[22] = N1042;
  assign OUT2[23] = N1043;
  assign OUT2[24] = N1044;
  assign OUT2[25] = N1045;
  assign OUT2[26] = N1046;
  assign OUT2[27] = N1047;
  assign OUT2[28] = N1048;
  assign OUT2[29] = N1049;
  assign OUT2[30] = N1050;
  assign OUT2[31] = N1051;

  AND3_X2 U1686 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .A3(RD1), .ZN(n1460) );
  AND3_X2 U1699 ( .A1(ADD_RD1[3]), .A2(n10665), .A3(RD1), .ZN(n1470) );
  AND3_X2 U1716 ( .A1(ADD_RD1[4]), .A2(n10658), .A3(RD1), .ZN(n1458) );
  AND3_X2 U1722 ( .A1(n10658), .A2(n10665), .A3(RD1), .ZN(n1477) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(n3005), .CK(CLK), .RN(n9883), .Q(n10538), .QN(n2102) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(n3004), .CK(CLK), .RN(n9883), .Q(n10539), .QN(n2110) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(n3003), .CK(CLK), .RN(n9883), .Q(n10540), .QN(n2118) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(n3002), .CK(CLK), .RN(n9883), .Q(n10541), .QN(n2126) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(n3001), .CK(CLK), .RN(n9883), .Q(n10542), .QN(n2134) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(n3000), .CK(CLK), .RN(n9883), .Q(n10543), .QN(n2142) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(n2999), .CK(CLK), .RN(n9883), .Q(n10544), .QN(n2150) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(n2998), .CK(CLK), .RN(n9883), .Q(n10545), .QN(n2158) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(n3133), .CK(CLK), .RN(n9883), .Q(n10562), .QN(n8326) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(n3132), .CK(CLK), .RN(n9883), .Q(n10563), .QN(n8325) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(n3131), .CK(CLK), .RN(n9883), .Q(n10564), .QN(n8324) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(n3130), .CK(CLK), .RN(n9883), .Q(n10565), .QN(n8323) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(n3129), .CK(CLK), .RN(n9883), .Q(n10566), .QN(n8322) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(n3128), .CK(CLK), .RN(n9883), .Q(n10567), .QN(n8321) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(n3127), .CK(CLK), .RN(n9883), .Q(n10568), .QN(n8320) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(n3126), .CK(CLK), .RN(n9883), .Q(n10569), .QN(n8319) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(n2973), .CK(CLK), .RN(n9883), .Q(n10554), .QN(n8342) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(n2972), .CK(CLK), .RN(n9883), .Q(n10555), .QN(n8341) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(n2971), .CK(CLK), .RN(n9883), .Q(n10556), .QN(n8340) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(n2970), .CK(CLK), .RN(n9883), .Q(n10557), .QN(n8339) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(n2969), .CK(CLK), .RN(n9883), .Q(n10558), .QN(n8338) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(n2968), .CK(CLK), .RN(n9883), .Q(n10559), .QN(n8337) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(n2967), .CK(CLK), .RN(n9883), .Q(n10560), .QN(n8336) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(n2966), .CK(CLK), .RN(n9883), .Q(n10561), .QN(n8335) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(n3101), .CK(CLK), .RN(n9883), .QN(n8509) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(n3100), .CK(CLK), .RN(n9883), .QN(n8508) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(n3099), .CK(CLK), .RN(n9883), .QN(n8507) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(n3098), .CK(CLK), .RN(n9883), .QN(n8506) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(n3097), .CK(CLK), .RN(n9883), .QN(n8505) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(n3096), .CK(CLK), .RN(n9883), .QN(n8504) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(n3095), .CK(CLK), .RN(n9883), .QN(n8503) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(n3094), .CK(CLK), .RN(n9883), .QN(n8502) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(n3069), .CK(CLK), .RN(n9883), .QN(n8334) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(n3068), .CK(CLK), .RN(n9883), .QN(n8333) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(n3067), .CK(CLK), .RN(n9883), .QN(n8332) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(n3066), .CK(CLK), .RN(n9883), .QN(n8331) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(n3065), .CK(CLK), .RN(n9883), .QN(n8330) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(n3064), .CK(CLK), .RN(n9883), .QN(n8329) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(n3063), .CK(CLK), .RN(n9883), .QN(n8328) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(n3062), .CK(CLK), .RN(n9883), .QN(n8327) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(n3165), .CK(CLK), .RN(n9883), .QN(n8597) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(n3164), .CK(CLK), .RN(n9883), .QN(n8596) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(n3163), .CK(CLK), .RN(n9883), .QN(n8595) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(n3162), .CK(CLK), .RN(n9883), .QN(n8594) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(n3161), .CK(CLK), .RN(n9883), .QN(n8593) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(n3160), .CK(CLK), .RN(n9883), .QN(n8592) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(n3159), .CK(CLK), .RN(n9883), .QN(n8591) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(n3158), .CK(CLK), .RN(n9883), .QN(n8590) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(n3811), .CK(CLK), .RN(n9883), .Q(n10432), 
        .QN(n8448) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(n9151), .CK(CLK), .RN(n9883), .Q(n10280), 
        .QN(n2276) );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(n9023), .CK(CLK), .RN(n9883), .Q(n10096), 
        .QN(n8227) );
  DFFR_X1 \REGISTERS_reg[0][9]  ( .D(n8959), .CK(CLK), .RN(n9883), .Q(n9944), 
        .QN(n2280) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(n9102), .CK(CLK), .RN(n9883), .Q(n10530), 
        .QN(n2295) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(n9103), .CK(CLK), .RN(n9883), .Q(n10531), 
        .QN(n2303) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(n9104), .CK(CLK), .RN(n9883), .Q(n10532), 
        .QN(n2311) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(n9105), .CK(CLK), .RN(n9883), .Q(n10533), 
        .QN(n2319) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(n9106), .CK(CLK), .RN(n9883), .Q(n10534), 
        .QN(n2327) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(n3846), .CK(CLK), .RN(n9883), .Q(n10498), 
        .QN(n8350) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(n3862), .CK(CLK), .RN(n9883), .Q(n10499), 
        .QN(n8349) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(n3878), .CK(CLK), .RN(n9883), .Q(n10500), 
        .QN(n8348) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(n3894), .CK(CLK), .RN(n9883), .Q(n10501), 
        .QN(n8347) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(n3910), .CK(CLK), .RN(n9883), .Q(n10502), 
        .QN(n8346) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(n3845), .CK(CLK), .RN(n9883), .QN(n8382)
         );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(n3861), .CK(CLK), .RN(n9883), .QN(n8381)
         );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(n3877), .CK(CLK), .RN(n9883), .QN(n8380)
         );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(n3893), .CK(CLK), .RN(n9883), .QN(n8379)
         );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(n3909), .CK(CLK), .RN(n9883), .QN(n8378)
         );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(n9134), .CK(CLK), .RN(n9883), .Q(n10626), 
        .QN(n8230) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(n9135), .CK(CLK), .RN(n9883), .Q(n10627), 
        .QN(n8232) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(n9136), .CK(CLK), .RN(n9883), .Q(n10628), 
        .QN(n8234) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(n9137), .CK(CLK), .RN(n9883), .Q(n10629), 
        .QN(n8236) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(n9138), .CK(CLK), .RN(n9883), .Q(n10630), 
        .QN(n8238) );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(n3844), .CK(CLK), .RN(n9883), .Q(n10466), 
        .QN(n8414) );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(n3860), .CK(CLK), .RN(n9883), .Q(n10467), 
        .QN(n8413) );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(n3876), .CK(CLK), .RN(n9883), .Q(n10468), 
        .QN(n8412) );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(n3892), .CK(CLK), .RN(n9883), .Q(n10469), 
        .QN(n8411) );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(n3908), .CK(CLK), .RN(n9883), .Q(n10470), 
        .QN(n8410) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(n3459), .CK(CLK), .RN(n9883), .Q(n10410), .QN(n8470) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(n3827), .CK(CLK), .RN(n9883), .Q(n10433), 
        .QN(n8447) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(n3843), .CK(CLK), .RN(n9883), .Q(n10434), 
        .QN(n8446) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(n3859), .CK(CLK), .RN(n9883), .Q(n10435), 
        .QN(n8445) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(n3875), .CK(CLK), .RN(n9883), .Q(n10436), 
        .QN(n8444) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(n3891), .CK(CLK), .RN(n9883), .Q(n10437), 
        .QN(n8443) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(n3907), .CK(CLK), .RN(n9883), .Q(n10438), 
        .QN(n8442) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(n3842), .CK(CLK), .RN(n9883), .Q(n10402), 
        .QN(n8517) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(n3858), .CK(CLK), .RN(n9883), .Q(n10403), 
        .QN(n8516) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(n3874), .CK(CLK), .RN(n9883), .Q(n10404), 
        .QN(n8515) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(n3890), .CK(CLK), .RN(n9883), .Q(n10405), 
        .QN(n8514) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(n3906), .CK(CLK), .RN(n9883), .Q(n10406), 
        .QN(n8513) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(n9173), .CK(CLK), .RN(n9883), .Q(n10258), .QN(n2100) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(n9150), .CK(CLK), .RN(n9883), .Q(n10281), 
        .QN(n2284) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(n9149), .CK(CLK), .RN(n9883), .Q(n10282), 
        .QN(n2292) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(n9148), .CK(CLK), .RN(n9883), .Q(n10283), 
        .QN(n2300) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(n9147), .CK(CLK), .RN(n9883), .Q(n10284), 
        .QN(n2308) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(n9146), .CK(CLK), .RN(n9883), .Q(n10285), 
        .QN(n2316) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(n9145), .CK(CLK), .RN(n9883), .Q(n10286), 
        .QN(n2324) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(n9077), .CK(CLK), .RN(n9883), .Q(n10226), .QN(n2107) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(n9045), .CK(CLK), .RN(n9883), .Q(n10074), 
        .QN(n8183) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(n9022), .CK(CLK), .RN(n9883), .Q(n10097), 
        .QN(n8229) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(n9021), .CK(CLK), .RN(n9883), .Q(n10098), 
        .QN(n8231) );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(n9020), .CK(CLK), .RN(n9883), .Q(n10099), 
        .QN(n8233) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(n9019), .CK(CLK), .RN(n9883), .Q(n10100), 
        .QN(n8235) );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(n9018), .CK(CLK), .RN(n9883), .Q(n10101), 
        .QN(n8237) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(n9017), .CK(CLK), .RN(n9883), .Q(n10102), 
        .QN(n8239) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(n9013), .CK(CLK), .RN(n9883), .Q(n10010), 
        .QN(n2105) );
  DFFR_X1 \REGISTERS_reg[0][31]  ( .D(n8981), .CK(CLK), .RN(n9883), .Q(n9922), 
        .QN(n2104) );
  DFFR_X1 \REGISTERS_reg[0][8]  ( .D(n8958), .CK(CLK), .RN(n9883), .Q(n9945), 
        .QN(n2288) );
  DFFR_X1 \REGISTERS_reg[0][7]  ( .D(n8957), .CK(CLK), .RN(n9883), .Q(n9946), 
        .QN(n2296) );
  DFFR_X1 \REGISTERS_reg[0][6]  ( .D(n8956), .CK(CLK), .RN(n9883), .Q(n9947), 
        .QN(n2304) );
  DFFR_X1 \REGISTERS_reg[0][5]  ( .D(n8955), .CK(CLK), .RN(n9883), .Q(n9948), 
        .QN(n2312) );
  DFFR_X1 \REGISTERS_reg[0][4]  ( .D(n8954), .CK(CLK), .RN(n9883), .Q(n9949), 
        .QN(n2320) );
  DFFR_X1 \REGISTERS_reg[0][3]  ( .D(n8953), .CK(CLK), .RN(n9883), .Q(n9950), 
        .QN(n2328) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(n3840), .CK(CLK), .RN(n9883), .Q(n10314), 
        .QN(n8605) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(n3856), .CK(CLK), .RN(n9883), .Q(n10315), 
        .QN(n8604) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(n3872), .CK(CLK), .RN(n9883), .Q(n10316), 
        .QN(n8603) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(n3888), .CK(CLK), .RN(n9883), .Q(n10317), 
        .QN(n8602) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(n3904), .CK(CLK), .RN(n9883), .Q(n10318), 
        .QN(n8601) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(n3197), .CK(CLK), .RN(n9883), .QN(n8302) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(n3229), .CK(CLK), .RN(n9883), .QN(n8685) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(n3837), .CK(CLK), .RN(n9883), .Q(n10218), 
        .QN(n8693) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(n3853), .CK(CLK), .RN(n9883), .Q(n10219), 
        .QN(n8692) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(n3869), .CK(CLK), .RN(n9883), .Q(n10220), 
        .QN(n8691) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(n3885), .CK(CLK), .RN(n9883), .Q(n10221), 
        .QN(n8690) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(n3901), .CK(CLK), .RN(n9883), .Q(n10222), 
        .QN(n8689) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(n3261), .CK(CLK), .RN(n9883), .Q(n10578), .QN(n8294) );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(n3293), .CK(CLK), .RN(n9883), .Q(n10138), .QN(n8773) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(n3836), .CK(CLK), .RN(n9883), .Q(n10130), 
        .QN(n2298) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(n3852), .CK(CLK), .RN(n9883), .Q(n10131), 
        .QN(n2306) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(n3868), .CK(CLK), .RN(n9883), .Q(n10132), 
        .QN(n2314) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(n3884), .CK(CLK), .RN(n9883), .Q(n10133), 
        .QN(n2322) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(n3900), .CK(CLK), .RN(n9883), .Q(n10134), 
        .QN(n2330) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(n3325), .CK(CLK), .RN(n9883), .QN(n8318)
         );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(n3357), .CK(CLK), .RN(n9883), .QN(n8829)
         );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(n3834), .CK(CLK), .RN(n9883), .Q(n10066), 
        .QN(n8837) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(n3850), .CK(CLK), .RN(n9883), .Q(n10067), 
        .QN(n8836) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(n3866), .CK(CLK), .RN(n9883), .Q(n10068), 
        .QN(n8835) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(n3882), .CK(CLK), .RN(n9883), .Q(n10069), 
        .QN(n8834) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(n3898), .CK(CLK), .RN(n9883), .Q(n10070), 
        .QN(n8833) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(n3389), .CK(CLK), .RN(n9883), .Q(n10570), 
        .QN(n8310) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(n3421), .CK(CLK), .RN(n9883), .QN(n8917)
         );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(n3832), .CK(CLK), .RN(n9883), .Q(n9978), 
        .QN(n8925) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(n3848), .CK(CLK), .RN(n9883), .Q(n9979), 
        .QN(n8924) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(n3864), .CK(CLK), .RN(n9883), .Q(n9980), 
        .QN(n8923) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(n3880), .CK(CLK), .RN(n9883), .Q(n9981), 
        .QN(n8922) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(n3896), .CK(CLK), .RN(n9883), .Q(n9982), 
        .QN(n8921) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(n3175), .CK(CLK), .RN(n9883), .QN(n8639)
         );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(n3174), .CK(CLK), .RN(n9883), .QN(n8638)
         );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(n3173), .CK(CLK), .RN(n9883), .QN(n8637)
         );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(n3172), .CK(CLK), .RN(n9883), .QN(n8636)
         );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(n3171), .CK(CLK), .RN(n9883), .QN(n8635)
         );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(n3170), .CK(CLK), .RN(n9883), .QN(n8634)
         );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(n3169), .CK(CLK), .RN(n9883), .QN(n8633)
         );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(n9055), .CK(CLK), .RN(n9883), .Q(n10248), 
        .QN(n2283) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(n9054), .CK(CLK), .RN(n9883), .Q(n10249), 
        .QN(n2291) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(n9053), .CK(CLK), .RN(n9883), .Q(n10250), 
        .QN(n2299) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(n9052), .CK(CLK), .RN(n9883), .Q(n10251), 
        .QN(n2307) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(n9051), .CK(CLK), .RN(n9883), .Q(n10252), 
        .QN(n2315) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(n9050), .CK(CLK), .RN(n9883), .Q(n10253), 
        .QN(n2323) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(n9049), .CK(CLK), .RN(n9883), .Q(n10254), 
        .QN(n2331) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(n3303), .CK(CLK), .RN(n9883), .QN(n8783)
         );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(n3302), .CK(CLK), .RN(n9883), .QN(n8782)
         );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(n3301), .CK(CLK), .RN(n9883), .QN(n8781)
         );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(n3300), .CK(CLK), .RN(n9883), .QN(n8780)
         );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(n3299), .CK(CLK), .RN(n9883), .QN(n8779)
         );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(n3298), .CK(CLK), .RN(n9883), .QN(n8778)
         );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(n3297), .CK(CLK), .RN(n9883), .QN(n8777)
         );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(n3450), .CK(CLK), .RN(n9883), .Q(n10042), 
        .QN(n8861) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(n3802), .CK(CLK), .RN(n9883), .Q(n10064), 
        .QN(n8839) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(n3818), .CK(CLK), .RN(n9883), .Q(n10065), 
        .QN(n8838) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(n9110), .CK(CLK), .RN(n9883), .Q(n10546), .QN(n8182) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(n9132), .CK(CLK), .RN(n9883), .Q(n10624), 
        .QN(n8226) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(n9133), .CK(CLK), .RN(n9883), .Q(n10625), 
        .QN(n8228) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(n3271), .CK(CLK), .RN(n9883), .Q(n10160), 
        .QN(n8751) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(n3270), .CK(CLK), .RN(n9883), .Q(n10161), 
        .QN(n8750) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(n3269), .CK(CLK), .RN(n9883), .Q(n10162), 
        .QN(n8749) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(n3268), .CK(CLK), .RN(n9883), .Q(n10163), 
        .QN(n8748) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(n3267), .CK(CLK), .RN(n9883), .Q(n10164), 
        .QN(n8747) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(n3266), .CK(CLK), .RN(n9883), .Q(n10165), 
        .QN(n8746) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(n3265), .CK(CLK), .RN(n9883), .Q(n10166), 
        .QN(n8745) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(n3399), .CK(CLK), .RN(n9883), .QN(n8895)
         );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(n3398), .CK(CLK), .RN(n9883), .QN(n8894)
         );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(n3397), .CK(CLK), .RN(n9883), .QN(n8893)
         );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(n3396), .CK(CLK), .RN(n9883), .QN(n8892)
         );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(n3395), .CK(CLK), .RN(n9883), .QN(n8891)
         );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(n3394), .CK(CLK), .RN(n9883), .QN(n8890)
         );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(n3393), .CK(CLK), .RN(n9883), .QN(n8889)
         );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(n3461), .CK(CLK), .RN(n9883), .QN(n8406) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(n3813), .CK(CLK), .RN(n9883), .QN(n8384)
         );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(n3829), .CK(CLK), .RN(n9883), .QN(n8383)
         );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(n3453), .CK(CLK), .RN(n9883), .Q(n10194), .QN(n8717) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(n3805), .CK(CLK), .RN(n9883), .Q(n10216), 
        .QN(n8695) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(n3821), .CK(CLK), .RN(n9883), .Q(n10217), 
        .QN(n8694) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(n8991), .CK(CLK), .RN(n9883), .Q(n10032), 
        .QN(n2281) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(n8990), .CK(CLK), .RN(n9883), .Q(n10033), 
        .QN(n2289) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(n8989), .CK(CLK), .RN(n9883), .Q(n10034), 
        .QN(n2297) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(n8988), .CK(CLK), .RN(n9883), .Q(n10035), 
        .QN(n2305) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(n8987), .CK(CLK), .RN(n9883), .Q(n10036), 
        .QN(n2313) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(n8986), .CK(CLK), .RN(n9883), .Q(n10037), 
        .QN(n2321) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(n8985), .CK(CLK), .RN(n9883), .Q(n10038), 
        .QN(n2329) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(n2997), .CK(CLK), .RN(n9883), .Q(n10586), .QN(n2166) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(n2996), .CK(CLK), .RN(n9883), .Q(n10587), .QN(n2174) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(n2995), .CK(CLK), .RN(n9883), .Q(n10588), .QN(n2182) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(n2994), .CK(CLK), .RN(n9883), .Q(n10589), .QN(n2190) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(n2993), .CK(CLK), .RN(n9883), .Q(n10590), .QN(n2198) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(n2992), .CK(CLK), .RN(n9883), .Q(n10591), .QN(n2206) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(n2991), .CK(CLK), .RN(n9883), .Q(n10592), .QN(n2214) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(n2990), .CK(CLK), .RN(n9883), .Q(n10593), .QN(n2222) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(n2989), .CK(CLK), .RN(n9883), .Q(n10594), .QN(n2230) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(n2988), .CK(CLK), .RN(n9883), .Q(n10595), .QN(n2238) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(n2987), .CK(CLK), .RN(n9883), .Q(n10596), .QN(n2246) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(n2986), .CK(CLK), .RN(n9883), .Q(n10597), .QN(n2254) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(n2985), .CK(CLK), .RN(n9883), .Q(n10598), .QN(n2262) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(n2984), .CK(CLK), .RN(n9883), .Q(n10599), .QN(n2270) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(n2983), .CK(CLK), .RN(n9883), .Q(n10600), 
        .QN(n2278) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(n2982), .CK(CLK), .RN(n9883), .Q(n10601), 
        .QN(n2286) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(n2981), .CK(CLK), .RN(n9883), .Q(n10602), 
        .QN(n2294) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(n2980), .CK(CLK), .RN(n9883), .Q(n10603), 
        .QN(n2302) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(n2979), .CK(CLK), .RN(n9883), .Q(n10604), 
        .QN(n2310) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(n2978), .CK(CLK), .RN(n9883), .Q(n10605), 
        .QN(n2318) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(n2977), .CK(CLK), .RN(n9883), .Q(n10606), 
        .QN(n2326) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(n2976), .CK(CLK), .RN(n9883), .Q(n10607), 
        .QN(n2334) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(n2975), .CK(CLK), .RN(n9883), .Q(n10608), 
        .QN(n2342) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(n2974), .CK(CLK), .RN(n9883), .Q(n10609), 
        .QN(n2350) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(n3460), .CK(CLK), .RN(n9883), .Q(n10442), .QN(n8438) );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(n3812), .CK(CLK), .RN(n9883), .Q(n10464), 
        .QN(n8416) );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(n3828), .CK(CLK), .RN(n9883), .Q(n10465), 
        .QN(n8415) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(n3125), .CK(CLK), .RN(n9883), .Q(n10322), .QN(n8565) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(n3124), .CK(CLK), .RN(n9883), .Q(n10323), .QN(n8564) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(n3123), .CK(CLK), .RN(n9883), .Q(n10324), .QN(n8563) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(n3122), .CK(CLK), .RN(n9883), .Q(n10325), .QN(n8562) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(n3121), .CK(CLK), .RN(n9883), .Q(n10326), .QN(n8561) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(n3120), .CK(CLK), .RN(n9883), .Q(n10327), .QN(n8560) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(n3119), .CK(CLK), .RN(n9883), .Q(n10328), .QN(n8559) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(n3118), .CK(CLK), .RN(n9883), .Q(n10329), .QN(n8558) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(n3117), .CK(CLK), .RN(n9883), .Q(n10330), .QN(n8557) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(n3116), .CK(CLK), .RN(n9883), .Q(n10331), .QN(n8556) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(n3115), .CK(CLK), .RN(n9883), .Q(n10332), .QN(n8555) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(n3114), .CK(CLK), .RN(n9883), .Q(n10333), .QN(n8554) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(n3113), .CK(CLK), .RN(n9883), .Q(n10334), .QN(n8553) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(n3112), .CK(CLK), .RN(n9883), .Q(n10335), .QN(n8552) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(n3111), .CK(CLK), .RN(n9883), .Q(n10336), 
        .QN(n8551) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(n3110), .CK(CLK), .RN(n9883), .Q(n10337), 
        .QN(n8550) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(n3109), .CK(CLK), .RN(n9883), .Q(n10338), 
        .QN(n8549) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(n3108), .CK(CLK), .RN(n9883), .Q(n10339), 
        .QN(n8548) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(n3107), .CK(CLK), .RN(n9883), .Q(n10340), 
        .QN(n8547) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(n3106), .CK(CLK), .RN(n9883), .Q(n10341), 
        .QN(n8546) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(n3105), .CK(CLK), .RN(n9883), .Q(n10342), 
        .QN(n8545) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(n3104), .CK(CLK), .RN(n9883), .Q(n10343), 
        .QN(n8544) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(n3103), .CK(CLK), .RN(n9883), .Q(n10344), 
        .QN(n8543) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(n3102), .CK(CLK), .RN(n9883), .Q(n10345), 
        .QN(n8542) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(n3456), .CK(CLK), .RN(n9883), .Q(n10290), .QN(n8629) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(n3808), .CK(CLK), .RN(n9883), .Q(n10312), 
        .QN(n8607) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(n3824), .CK(CLK), .RN(n9883), .Q(n10313), 
        .QN(n8606) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(n3239), .CK(CLK), .RN(n9883), .Q(n10184), 
        .QN(n8727) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(n3238), .CK(CLK), .RN(n9883), .Q(n10185), 
        .QN(n8726) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(n3237), .CK(CLK), .RN(n9883), .Q(n10186), 
        .QN(n8725) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(n3236), .CK(CLK), .RN(n9883), .Q(n10187), 
        .QN(n8724) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(n3235), .CK(CLK), .RN(n9883), .Q(n10188), 
        .QN(n8723) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(n3234), .CK(CLK), .RN(n9883), .Q(n10189), 
        .QN(n8722) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(n3233), .CK(CLK), .RN(n9883), .Q(n10190), 
        .QN(n8721) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(n3452), .CK(CLK), .RN(n9883), .Q(n10106), 
        .QN(n2106) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(n3804), .CK(CLK), .RN(n9883), .Q(n10128), 
        .QN(n2282) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(n3820), .CK(CLK), .RN(n9883), .Q(n10129), 
        .QN(n2290) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(n3367), .CK(CLK), .RN(n9883), .Q(n10000), 
        .QN(n8871) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(n3366), .CK(CLK), .RN(n9883), .Q(n10001), 
        .QN(n8870) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(n3365), .CK(CLK), .RN(n9883), .Q(n10002), 
        .QN(n8869) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(n3364), .CK(CLK), .RN(n9883), .Q(n10003), 
        .QN(n8868) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(n3363), .CK(CLK), .RN(n9883), .Q(n10004), 
        .QN(n8867) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(n3362), .CK(CLK), .RN(n9883), .Q(n10005), 
        .QN(n8866) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(n3361), .CK(CLK), .RN(n9883), .Q(n10006), 
        .QN(n8865) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(n3448), .CK(CLK), .RN(n9883), .Q(n9954), 
        .QN(n8949) );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(n3800), .CK(CLK), .RN(n9883), .Q(n9976), 
        .QN(n8927) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(n3816), .CK(CLK), .RN(n9883), .Q(n9977), 
        .QN(n8926) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(n2965), .CK(CLK), .RN(n9883), .Q(n10634), .QN(n8286) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(n2964), .CK(CLK), .RN(n9883), .Q(n10635), .QN(n8285) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(n2963), .CK(CLK), .RN(n9883), .Q(n10636), .QN(n8284) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(n2962), .CK(CLK), .RN(n9883), .Q(n10637), .QN(n8283) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(n2961), .CK(CLK), .RN(n9883), .Q(n10638), .QN(n8282) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(n2960), .CK(CLK), .RN(n9883), .Q(n10639), .QN(n8281) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(n2959), .CK(CLK), .RN(n9883), .Q(n10640), .QN(n8280) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(n2958), .CK(CLK), .RN(n9883), .Q(n10641), .QN(n8279) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(n2957), .CK(CLK), .RN(n9883), .Q(n10642), .QN(n8278) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(n2956), .CK(CLK), .RN(n9883), .Q(n10643), .QN(n8277) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(n2955), .CK(CLK), .RN(n9883), .Q(n10644), .QN(n8276) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(n2954), .CK(CLK), .RN(n9883), .Q(n10645), .QN(n8275) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(n2953), .CK(CLK), .RN(n9883), .Q(n10646), .QN(n8274) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(n2952), .CK(CLK), .RN(n9883), .Q(n10647), .QN(n8273) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(n2951), .CK(CLK), .RN(n9883), .Q(n10648), 
        .QN(n8272) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(n2950), .CK(CLK), .RN(n9883), .Q(n10649), 
        .QN(n8271) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(n2949), .CK(CLK), .RN(n9883), .Q(n10650), 
        .QN(n8270) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(n2948), .CK(CLK), .RN(n9883), .Q(n10651), 
        .QN(n8269) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(n2947), .CK(CLK), .RN(n9883), .Q(n10652), 
        .QN(n8268) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(n2946), .CK(CLK), .RN(n9883), .Q(n10653), 
        .QN(n8267) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(n2945), .CK(CLK), .RN(n9883), .Q(n10654), 
        .QN(n8266) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(n2944), .CK(CLK), .RN(n9883), .Q(n10655), 
        .QN(n8265) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(n2943), .CK(CLK), .RN(n9883), .Q(n10656), 
        .QN(n8264) );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(n2942), .CK(CLK), .RN(n9883), .Q(n10657), 
        .QN(n8263) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(n3093), .CK(CLK), .RN(n9883), .QN(n8501) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(n3092), .CK(CLK), .RN(n9883), .QN(n8500) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(n3091), .CK(CLK), .RN(n9883), .QN(n8499) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(n3090), .CK(CLK), .RN(n9883), .QN(n8498) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(n3089), .CK(CLK), .RN(n9883), .QN(n8497) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(n3088), .CK(CLK), .RN(n9883), .QN(n8496) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(n3087), .CK(CLK), .RN(n9883), .QN(n8495) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(n3086), .CK(CLK), .RN(n9883), .QN(n8494) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(n3085), .CK(CLK), .RN(n9883), .QN(n8493) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(n3084), .CK(CLK), .RN(n9883), .QN(n8492) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(n3083), .CK(CLK), .RN(n9883), .QN(n8491) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(n3082), .CK(CLK), .RN(n9883), .QN(n8490) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(n3081), .CK(CLK), .RN(n9883), .QN(n8489) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(n3080), .CK(CLK), .RN(n9883), .QN(n8488) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(n3079), .CK(CLK), .RN(n9883), .QN(n8487)
         );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(n3078), .CK(CLK), .RN(n9883), .QN(n8486)
         );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(n3077), .CK(CLK), .RN(n9883), .QN(n8485)
         );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(n3076), .CK(CLK), .RN(n9883), .QN(n8484)
         );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(n3075), .CK(CLK), .RN(n9883), .QN(n8483)
         );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(n3074), .CK(CLK), .RN(n9883), .QN(n8482)
         );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(n3073), .CK(CLK), .RN(n9883), .QN(n8481)
         );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(n3072), .CK(CLK), .RN(n9883), .QN(n8480)
         );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(n3071), .CK(CLK), .RN(n9883), .QN(n8479)
         );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(n3070), .CK(CLK), .RN(n9883), .QN(n8478)
         );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(n3207), .CK(CLK), .RN(n9883), .QN(n8663)
         );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(n3206), .CK(CLK), .RN(n9883), .QN(n8662)
         );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(n3205), .CK(CLK), .RN(n9883), .QN(n8661)
         );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(n3204), .CK(CLK), .RN(n9883), .QN(n8660)
         );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(n3203), .CK(CLK), .RN(n9883), .QN(n8659)
         );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(n3202), .CK(CLK), .RN(n9883), .QN(n8658)
         );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(n3201), .CK(CLK), .RN(n9883), .QN(n8657)
         );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(n3335), .CK(CLK), .RN(n9883), .QN(n8807)
         );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(n3334), .CK(CLK), .RN(n9883), .QN(n8806)
         );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(n3333), .CK(CLK), .RN(n9883), .QN(n8805)
         );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(n3332), .CK(CLK), .RN(n9883), .QN(n8804)
         );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(n3331), .CK(CLK), .RN(n9883), .QN(n8803)
         );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(n3330), .CK(CLK), .RN(n9883), .QN(n8802)
         );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(n3329), .CK(CLK), .RN(n9883), .QN(n8801)
         );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(n9078), .CK(CLK), .RN(n9883), .Q(n10506), .QN(n2103) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(n9100), .CK(CLK), .RN(n9883), .Q(n10528), 
        .QN(n2279) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(n9101), .CK(CLK), .RN(n9883), .Q(n10529), 
        .QN(n2287) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(n3061), .CK(CLK), .RN(n9883), .QN(n8262) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(n3060), .CK(CLK), .RN(n9883), .QN(n8261) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(n3059), .CK(CLK), .RN(n9883), .QN(n8260) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(n3058), .CK(CLK), .RN(n9883), .QN(n8259) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(n3057), .CK(CLK), .RN(n9883), .QN(n8258) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(n3056), .CK(CLK), .RN(n9883), .QN(n8257) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(n3055), .CK(CLK), .RN(n9883), .QN(n8256) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(n3054), .CK(CLK), .RN(n9883), .QN(n8255) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(n3053), .CK(CLK), .RN(n9883), .QN(n8254) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(n3052), .CK(CLK), .RN(n9883), .QN(n8253) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(n3051), .CK(CLK), .RN(n9883), .QN(n8252) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(n3050), .CK(CLK), .RN(n9883), .QN(n8251) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(n3049), .CK(CLK), .RN(n9883), .QN(n8250) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(n3048), .CK(CLK), .RN(n9883), .QN(n8249) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(n3047), .CK(CLK), .RN(n9883), .QN(n8248)
         );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(n3046), .CK(CLK), .RN(n9883), .QN(n8247)
         );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(n3045), .CK(CLK), .RN(n9883), .QN(n8246)
         );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(n3044), .CK(CLK), .RN(n9883), .QN(n8477)
         );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(n3043), .CK(CLK), .RN(n9883), .QN(n8476)
         );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(n3042), .CK(CLK), .RN(n9883), .QN(n8475)
         );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(n3041), .CK(CLK), .RN(n9883), .QN(n8474)
         );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(n3040), .CK(CLK), .RN(n9883), .QN(n8473)
         );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(n3039), .CK(CLK), .RN(n9883), .QN(n8472)
         );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(n3038), .CK(CLK), .RN(n9883), .QN(n8471)
         );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(n3462), .CK(CLK), .RN(n9883), .Q(n10474), .QN(n8374) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(n3814), .CK(CLK), .RN(n9883), .Q(n10496), 
        .QN(n8352) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(n3830), .CK(CLK), .RN(n9883), .Q(n10497), 
        .QN(n8351) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(n3458), .CK(CLK), .RN(n9883), .Q(n10378), .QN(n8541) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(n3810), .CK(CLK), .RN(n9883), .Q(n10400), 
        .QN(n8519) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(n3826), .CK(CLK), .RN(n9883), .Q(n10401), 
        .QN(n8518) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(n9205), .CK(CLK), .RN(n9878), .Q(n10346), .QN(n2101) );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(n3157), .CK(CLK), .RN(n9883), .QN(n8589) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(n3156), .CK(CLK), .RN(n9883), .QN(n8588) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(n3155), .CK(CLK), .RN(n9883), .QN(n8587) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(n3154), .CK(CLK), .RN(n9883), .QN(n8586) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(n3153), .CK(CLK), .RN(n9883), .QN(n8585) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(n3152), .CK(CLK), .RN(n9883), .QN(n8584) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(n3151), .CK(CLK), .RN(n9883), .QN(n8583) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(n3150), .CK(CLK), .RN(n9883), .QN(n8582) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(n3149), .CK(CLK), .RN(n9883), .QN(n8581) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(n3148), .CK(CLK), .RN(n9883), .QN(n8580) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(n3147), .CK(CLK), .RN(n9883), .QN(n8579) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(n3146), .CK(CLK), .RN(n9883), .QN(n8578) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(n3145), .CK(CLK), .RN(n9883), .QN(n8577) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(n3144), .CK(CLK), .RN(n9883), .QN(n8576) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(n3143), .CK(CLK), .RN(n9883), .QN(n8575)
         );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(n3142), .CK(CLK), .RN(n9883), .QN(n8574)
         );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(n3141), .CK(CLK), .RN(n9883), .QN(n8573)
         );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(n3140), .CK(CLK), .RN(n9883), .QN(n8572)
         );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(n3139), .CK(CLK), .RN(n9883), .QN(n8571)
         );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(n3138), .CK(CLK), .RN(n9883), .QN(n8570)
         );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(n3137), .CK(CLK), .RN(n9883), .QN(n8569)
         );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(n3136), .CK(CLK), .RN(n9883), .QN(n8568)
         );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(n3135), .CK(CLK), .RN(n9883), .QN(n8567)
         );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(n3134), .CK(CLK), .RN(n9883), .QN(n8566)
         );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(n9079), .CK(CLK), .RN(n9883), .Q(n10507), .QN(n2111) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(n9080), .CK(CLK), .RN(n9883), .Q(n10508), .QN(n2119) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(n9081), .CK(CLK), .RN(n9883), .Q(n10509), .QN(n2127) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(n9082), .CK(CLK), .RN(n9883), .Q(n10510), .QN(n2135) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(n9083), .CK(CLK), .RN(n9883), .Q(n10511), .QN(n2143) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(n9084), .CK(CLK), .RN(n9883), .Q(n10512), .QN(n2151) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(n9085), .CK(CLK), .RN(n9883), .Q(n10513), .QN(n2159) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(n9086), .CK(CLK), .RN(n9883), .Q(n10514), .QN(n2167) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(n9087), .CK(CLK), .RN(n9883), .Q(n10515), .QN(n2175) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(n9088), .CK(CLK), .RN(n9883), .Q(n10516), .QN(n2183) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(n9089), .CK(CLK), .RN(n9883), .Q(n10517), .QN(n2191) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(n9090), .CK(CLK), .RN(n9883), .Q(n10518), .QN(n2199) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(n9091), .CK(CLK), .RN(n9883), .Q(n10519), .QN(n2207) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(n9092), .CK(CLK), .RN(n9883), .Q(n10520), .QN(n2215) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(n9093), .CK(CLK), .RN(n9883), .Q(n10521), .QN(n2223) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(n9094), .CK(CLK), .RN(n9883), .Q(n10522), .QN(n2231) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(n9095), .CK(CLK), .RN(n9883), .Q(n10523), .QN(n2239) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(n9096), .CK(CLK), .RN(n9883), .Q(n10524), .QN(n2247) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(n9097), .CK(CLK), .RN(n9883), .Q(n10525), .QN(n2255) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(n9098), .CK(CLK), .RN(n9883), .Q(n10526), .QN(n2263) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(n9099), .CK(CLK), .RN(n9883), .Q(n10527), .QN(n2271) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(n9107), .CK(CLK), .RN(n9883), .Q(n10535), 
        .QN(n2335) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(n9108), .CK(CLK), .RN(n9883), .Q(n10536), 
        .QN(n2343) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(n9109), .CK(CLK), .RN(n9883), .Q(n10537), 
        .QN(n2351) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(n3478), .CK(CLK), .RN(n9883), .Q(n10475), .QN(n8373) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(n3494), .CK(CLK), .RN(n9883), .Q(n10476), .QN(n8372) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(n3510), .CK(CLK), .RN(n9883), .Q(n10477), .QN(n8371) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(n3526), .CK(CLK), .RN(n9883), .Q(n10478), .QN(n8370) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(n3542), .CK(CLK), .RN(n9883), .Q(n10479), .QN(n8369) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(n3558), .CK(CLK), .RN(n9883), .Q(n10480), .QN(n8368) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(n3574), .CK(CLK), .RN(n9883), .Q(n10481), .QN(n8367) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(n3590), .CK(CLK), .RN(n9883), .Q(n10482), .QN(n8366) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(n3606), .CK(CLK), .RN(n9883), .Q(n10483), .QN(n8365) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(n3622), .CK(CLK), .RN(n9883), .Q(n10484), .QN(n8364) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(n3638), .CK(CLK), .RN(n9883), .Q(n10485), .QN(n8363) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(n3654), .CK(CLK), .RN(n9883), .Q(n10486), .QN(n8362) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(n3670), .CK(CLK), .RN(n9883), .Q(n10487), .QN(n8361) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(n3686), .CK(CLK), .RN(n9883), .Q(n10488), .QN(n8360) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(n3702), .CK(CLK), .RN(n9883), .Q(n10489), .QN(n8359) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(n3718), .CK(CLK), .RN(n9883), .Q(n10490), .QN(n8358) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(n3734), .CK(CLK), .RN(n9883), .Q(n10491), .QN(n8357) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(n3750), .CK(CLK), .RN(n9883), .Q(n10492), .QN(n8356) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(n3766), .CK(CLK), .RN(n9883), .Q(n10493), .QN(n8355) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(n3782), .CK(CLK), .RN(n9883), .Q(n10494), .QN(n8354) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(n3798), .CK(CLK), .RN(n9883), .Q(n10495), .QN(n8353) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(n3926), .CK(CLK), .RN(n9883), .Q(n10503), 
        .QN(n8345) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(n3942), .CK(CLK), .RN(n9879), .Q(n10504), 
        .QN(n8344) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(n3958), .CK(CLK), .RN(n9883), .Q(n10505), 
        .QN(n8343) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(n3477), .CK(CLK), .RN(n9883), .QN(n8405) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(n3493), .CK(CLK), .RN(n9883), .QN(n8404) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(n3509), .CK(CLK), .RN(n9883), .QN(n8403) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(n3525), .CK(CLK), .RN(n9883), .QN(n8402) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(n3541), .CK(CLK), .RN(n9883), .QN(n8401) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(n3557), .CK(CLK), .RN(n9883), .QN(n8400) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(n3573), .CK(CLK), .RN(n9883), .QN(n8399) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(n3589), .CK(CLK), .RN(n9883), .QN(n8398) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(n3605), .CK(CLK), .RN(n9883), .QN(n8397) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(n3621), .CK(CLK), .RN(n9883), .QN(n8396) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(n3637), .CK(CLK), .RN(n9883), .QN(n8395) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(n3653), .CK(CLK), .RN(n9883), .QN(n8394) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(n3669), .CK(CLK), .RN(n9883), .QN(n8393) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(n3685), .CK(CLK), .RN(n9883), .QN(n8392) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(n3701), .CK(CLK), .RN(n9883), .QN(n8391) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(n3717), .CK(CLK), .RN(n9883), .QN(n8390) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(n3733), .CK(CLK), .RN(n9883), .QN(n8389) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(n3749), .CK(CLK), .RN(n9883), .QN(n8388) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(n3765), .CK(CLK), .RN(n9883), .QN(n8387) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(n3781), .CK(CLK), .RN(n9883), .QN(n8386) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(n3797), .CK(CLK), .RN(n9883), .QN(n8385) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(n3925), .CK(CLK), .RN(n9883), .QN(n8377)
         );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(n3941), .CK(CLK), .RN(n9879), .QN(n8376)
         );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(n3957), .CK(CLK), .RN(n9883), .QN(n8375)
         );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(n9111), .CK(CLK), .RN(n9883), .Q(n10547), .QN(n8184) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(n9112), .CK(CLK), .RN(n9883), .Q(n10548), .QN(n8186) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(n9113), .CK(CLK), .RN(n9883), .Q(n10549), .QN(n8188) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(n9114), .CK(CLK), .RN(n9883), .Q(n10550), .QN(n8190) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(n9115), .CK(CLK), .RN(n9883), .Q(n10551), .QN(n8192) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(n9116), .CK(CLK), .RN(n9883), .Q(n10552), .QN(n8194) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(n9117), .CK(CLK), .RN(n9883), .Q(n10553), .QN(n8196) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(n9118), .CK(CLK), .RN(n9883), .Q(n10610), .QN(n8198) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(n9119), .CK(CLK), .RN(n9883), .Q(n10611), .QN(n8200) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(n9120), .CK(CLK), .RN(n9883), .Q(n10612), .QN(n8202) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(n9121), .CK(CLK), .RN(n9883), .Q(n10613), .QN(n8204) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(n9122), .CK(CLK), .RN(n9883), .Q(n10614), .QN(n8206) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(n9123), .CK(CLK), .RN(n9883), .Q(n10615), .QN(n8208) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(n9124), .CK(CLK), .RN(n9883), .Q(n10616), .QN(n8210) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(n9125), .CK(CLK), .RN(n9883), .Q(n10617), .QN(n8212) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(n9126), .CK(CLK), .RN(n9883), .Q(n10618), .QN(n8214) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(n9127), .CK(CLK), .RN(n9883), .Q(n10619), .QN(n8216) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(n9128), .CK(CLK), .RN(n9883), .Q(n10620), .QN(n8218) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(n9129), .CK(CLK), .RN(n9883), .Q(n10621), .QN(n8220) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(n9130), .CK(CLK), .RN(n9883), .Q(n10622), .QN(n8222) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(n9131), .CK(CLK), .RN(n9883), .Q(n10623), .QN(n8224) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(n9139), .CK(CLK), .RN(n9883), .Q(n10631), 
        .QN(n8240) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(n9140), .CK(CLK), .RN(n9883), .Q(n10632), 
        .QN(n8242) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(n9141), .CK(CLK), .RN(n9883), .Q(n10633), 
        .QN(n8244) );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(n3476), .CK(CLK), .RN(n9883), .Q(n10443), .QN(n8437) );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(n3492), .CK(CLK), .RN(n9883), .Q(n10444), .QN(n8436) );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(n3508), .CK(CLK), .RN(n9883), .Q(n10445), .QN(n8435) );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(n3524), .CK(CLK), .RN(n9883), .Q(n10446), .QN(n8434) );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(n3540), .CK(CLK), .RN(n9883), .Q(n10447), .QN(n8433) );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(n3556), .CK(CLK), .RN(n9883), .Q(n10448), .QN(n8432) );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(n3572), .CK(CLK), .RN(n9883), .Q(n10449), .QN(n8431) );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(n3588), .CK(CLK), .RN(n9883), .Q(n10450), .QN(n8430) );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(n3604), .CK(CLK), .RN(n9883), .Q(n10451), .QN(n8429) );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(n3620), .CK(CLK), .RN(n9883), .Q(n10452), .QN(n8428) );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(n3636), .CK(CLK), .RN(n9883), .Q(n10453), .QN(n8427) );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(n3652), .CK(CLK), .RN(n9883), .Q(n10454), .QN(n8426) );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(n3668), .CK(CLK), .RN(n9883), .Q(n10455), .QN(n8425) );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(n3684), .CK(CLK), .RN(n9883), .Q(n10456), .QN(n8424) );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(n3700), .CK(CLK), .RN(n9883), .Q(n10457), .QN(n8423) );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(n3716), .CK(CLK), .RN(n9883), .Q(n10458), .QN(n8422) );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(n3732), .CK(CLK), .RN(n9883), .Q(n10459), .QN(n8421) );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(n3748), .CK(CLK), .RN(n9883), .Q(n10460), .QN(n8420) );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(n3764), .CK(CLK), .RN(n9883), .Q(n10461), .QN(n8419) );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(n3780), .CK(CLK), .RN(n9883), .Q(n10462), .QN(n8418) );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(n3796), .CK(CLK), .RN(n9883), .Q(n10463), .QN(n8417) );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(n3924), .CK(CLK), .RN(n9883), .Q(n10471), 
        .QN(n8409) );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(n3940), .CK(CLK), .RN(n9879), .Q(n10472), 
        .QN(n8408) );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(n3956), .CK(CLK), .RN(n9883), .Q(n10473), 
        .QN(n8407) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(n3475), .CK(CLK), .RN(n9883), .Q(n10411), .QN(n8469) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(n3491), .CK(CLK), .RN(n9883), .Q(n10412), .QN(n8468) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(n3507), .CK(CLK), .RN(n9883), .Q(n10413), .QN(n8467) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(n3523), .CK(CLK), .RN(n9883), .Q(n10414), .QN(n8466) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(n3539), .CK(CLK), .RN(n9883), .Q(n10415), .QN(n8465) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(n3555), .CK(CLK), .RN(n9883), .Q(n10416), .QN(n8464) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(n3571), .CK(CLK), .RN(n9883), .Q(n10417), .QN(n8463) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(n3587), .CK(CLK), .RN(n9883), .Q(n10418), .QN(n8462) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(n3603), .CK(CLK), .RN(n9883), .Q(n10419), .QN(n8461) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(n3619), .CK(CLK), .RN(n9883), .Q(n10420), .QN(n8460) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(n3635), .CK(CLK), .RN(n9883), .Q(n10421), .QN(n8459) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(n3651), .CK(CLK), .RN(n9883), .Q(n10422), .QN(n8458) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(n3667), .CK(CLK), .RN(n9883), .Q(n10423), .QN(n8457) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(n3683), .CK(CLK), .RN(n9883), .Q(n10424), .QN(n8456) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(n3699), .CK(CLK), .RN(n9883), .Q(n10425), .QN(n8455) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(n3715), .CK(CLK), .RN(n9883), .Q(n10426), .QN(n8454) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(n3731), .CK(CLK), .RN(n9883), .Q(n10427), .QN(n8453) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(n3747), .CK(CLK), .RN(n9883), .Q(n10428), .QN(n8452) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(n3763), .CK(CLK), .RN(n9883), .Q(n10429), .QN(n8451) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(n3779), .CK(CLK), .RN(n9883), .Q(n10430), .QN(n8450) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(n3795), .CK(CLK), .RN(n9883), .Q(n10431), .QN(n8449) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(n3923), .CK(CLK), .RN(n9883), .Q(n10439), 
        .QN(n8441) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(n3939), .CK(CLK), .RN(n9879), .Q(n10440), 
        .QN(n8440) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(n3955), .CK(CLK), .RN(n9883), .Q(n10441), 
        .QN(n8439) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(n3474), .CK(CLK), .RN(n9883), .Q(n10379), .QN(n8540) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(n3490), .CK(CLK), .RN(n9883), .Q(n10380), .QN(n8539) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(n3506), .CK(CLK), .RN(n9883), .Q(n10381), .QN(n8538) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(n3522), .CK(CLK), .RN(n9883), .Q(n10382), .QN(n8537) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(n3538), .CK(CLK), .RN(n9883), .Q(n10383), .QN(n8536) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(n3554), .CK(CLK), .RN(n9883), .Q(n10384), .QN(n8535) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(n3570), .CK(CLK), .RN(n9883), .Q(n10385), .QN(n8534) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(n3586), .CK(CLK), .RN(n9883), .Q(n10386), .QN(n8533) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(n3602), .CK(CLK), .RN(n9883), .Q(n10387), .QN(n8532) );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(n3618), .CK(CLK), .RN(n9883), .Q(n10388), .QN(n8531) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(n3634), .CK(CLK), .RN(n9883), .Q(n10389), .QN(n8530) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(n3650), .CK(CLK), .RN(n9883), .Q(n10390), .QN(n8529) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(n3666), .CK(CLK), .RN(n9883), .Q(n10391), .QN(n8528) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(n3682), .CK(CLK), .RN(n9883), .Q(n10392), .QN(n8527) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(n3698), .CK(CLK), .RN(n9883), .Q(n10393), .QN(n8526) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(n3714), .CK(CLK), .RN(n9883), .Q(n10394), .QN(n8525) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(n3730), .CK(CLK), .RN(n9883), .Q(n10395), .QN(n8524) );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(n3746), .CK(CLK), .RN(n9883), .Q(n10396), .QN(n8523) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(n3762), .CK(CLK), .RN(n9883), .Q(n10397), .QN(n8522) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(n3778), .CK(CLK), .RN(n9883), .Q(n10398), .QN(n8521) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(n3794), .CK(CLK), .RN(n9883), .Q(n10399), .QN(n8520) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(n3922), .CK(CLK), .RN(n9883), .Q(n10407), 
        .QN(n8512) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(n3938), .CK(CLK), .RN(n9883), .Q(n10408), 
        .QN(n8511) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(n3954), .CK(CLK), .RN(n9883), .Q(n10409), 
        .QN(n8510) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(n9172), .CK(CLK), .RN(n9883), .Q(n10259), .QN(n2108) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(n9171), .CK(CLK), .RN(n9883), .Q(n10260), .QN(n2116) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(n9170), .CK(CLK), .RN(n9883), .Q(n10261), .QN(n2124) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(n9169), .CK(CLK), .RN(n9883), .Q(n10262), .QN(n2132) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(n9168), .CK(CLK), .RN(n9883), .Q(n10263), .QN(n2140) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(n9167), .CK(CLK), .RN(n9883), .Q(n10264), .QN(n2148) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(n9166), .CK(CLK), .RN(n9883), .Q(n10265), .QN(n2156) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(n9165), .CK(CLK), .RN(n9883), .Q(n10266), .QN(n2164) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(n9164), .CK(CLK), .RN(n9883), .Q(n10267), .QN(n2172) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(n9163), .CK(CLK), .RN(n9883), .Q(n10268), .QN(n2180) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(n9162), .CK(CLK), .RN(n9883), .Q(n10269), .QN(n2188) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(n9161), .CK(CLK), .RN(n9883), .Q(n10270), .QN(n2196) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(n9160), .CK(CLK), .RN(n9883), .Q(n10271), .QN(n2204) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(n9159), .CK(CLK), .RN(n9883), .Q(n10272), .QN(n2212) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(n9158), .CK(CLK), .RN(n9883), .Q(n10273), .QN(n2220) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(n9157), .CK(CLK), .RN(n9883), .Q(n10274), .QN(n2228) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(n9156), .CK(CLK), .RN(n9883), .Q(n10275), .QN(n2236) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(n9155), .CK(CLK), .RN(n9883), .Q(n10276), .QN(n2244) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(n9154), .CK(CLK), .RN(n9883), .Q(n10277), .QN(n2252) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(n9153), .CK(CLK), .RN(n9883), .Q(n10278), .QN(n2260) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(n9152), .CK(CLK), .RN(n9883), .Q(n10279), .QN(n2268) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(n9144), .CK(CLK), .RN(n9883), .Q(n10287), 
        .QN(n2332) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(n9143), .CK(CLK), .RN(n9883), .Q(n10288), 
        .QN(n2340) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(n9142), .CK(CLK), .RN(n9883), .Q(n10289), 
        .QN(n2348) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(n9076), .CK(CLK), .RN(n9883), .Q(n10227), .QN(n2115) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(n9075), .CK(CLK), .RN(n9883), .Q(n10228), .QN(n2123) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(n9074), .CK(CLK), .RN(n9883), .Q(n10229), .QN(n2131) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(n9073), .CK(CLK), .RN(n9883), .Q(n10230), .QN(n2139) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(n9072), .CK(CLK), .RN(n9883), .Q(n10231), .QN(n2147) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(n9071), .CK(CLK), .RN(n9883), .Q(n10232), .QN(n2155) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(n9070), .CK(CLK), .RN(n9883), .Q(n10233), .QN(n2163) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(n9069), .CK(CLK), .RN(n9883), .Q(n10234), .QN(n2171) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(n9068), .CK(CLK), .RN(n9883), .Q(n10235), .QN(n2179) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(n9067), .CK(CLK), .RN(n9883), .Q(n10236), .QN(n2187) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(n9066), .CK(CLK), .RN(n9883), .Q(n10237), .QN(n2195) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(n9065), .CK(CLK), .RN(n9883), .Q(n10238), .QN(n2203) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(n9064), .CK(CLK), .RN(n9883), .Q(n10239), .QN(n2211) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(n9063), .CK(CLK), .RN(n9883), .Q(n10240), .QN(n2219) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(n9062), .CK(CLK), .RN(n9883), .Q(n10241), .QN(n2227) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(n9061), .CK(CLK), .RN(n9883), .Q(n10242), .QN(n2235) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(n9060), .CK(CLK), .RN(n9883), .Q(n10243), .QN(n2243) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(n9059), .CK(CLK), .RN(n9883), .Q(n10244), .QN(n2251) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(n9058), .CK(CLK), .RN(n9883), .Q(n10245), .QN(n2259) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(n9057), .CK(CLK), .RN(n9883), .Q(n10246), .QN(n2267) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(n9056), .CK(CLK), .RN(n9883), .Q(n10247), .QN(n2275) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(n9048), .CK(CLK), .RN(n9883), .Q(n10255), 
        .QN(n2339) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(n9047), .CK(CLK), .RN(n9883), .Q(n10256), 
        .QN(n2347) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(n9046), .CK(CLK), .RN(n9883), .Q(n10257), 
        .QN(n2355) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(n9044), .CK(CLK), .RN(n9883), .Q(n10075), 
        .QN(n8185) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(n9043), .CK(CLK), .RN(n9883), .Q(n10076), 
        .QN(n8187) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(n9042), .CK(CLK), .RN(n9883), .Q(n10077), 
        .QN(n8189) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(n9041), .CK(CLK), .RN(n9883), .Q(n10078), 
        .QN(n8191) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(n9040), .CK(CLK), .RN(n9883), .Q(n10079), 
        .QN(n8193) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(n9039), .CK(CLK), .RN(n9883), .Q(n10080), 
        .QN(n8195) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(n9038), .CK(CLK), .RN(n9883), .Q(n10081), 
        .QN(n8197) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(n9037), .CK(CLK), .RN(n9883), .Q(n10082), 
        .QN(n8199) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(n9036), .CK(CLK), .RN(n9883), .Q(n10083), 
        .QN(n8201) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(n9035), .CK(CLK), .RN(n9883), .Q(n10084), 
        .QN(n8203) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(n9034), .CK(CLK), .RN(n9883), .Q(n10085), 
        .QN(n8205) );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(n9033), .CK(CLK), .RN(n9883), .Q(n10086), 
        .QN(n8207) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(n9032), .CK(CLK), .RN(n9883), .Q(n10087), 
        .QN(n8209) );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(n9031), .CK(CLK), .RN(n9883), .Q(n10088), 
        .QN(n8211) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(n9030), .CK(CLK), .RN(n9883), .Q(n10089), 
        .QN(n8213) );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(n9029), .CK(CLK), .RN(n9883), .Q(n10090), 
        .QN(n8215) );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(n9028), .CK(CLK), .RN(n9883), .Q(n10091), 
        .QN(n8217) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(n9027), .CK(CLK), .RN(n9883), .Q(n10092), 
        .QN(n8219) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(n9026), .CK(CLK), .RN(n9883), .Q(n10093), 
        .QN(n8221) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(n9025), .CK(CLK), .RN(n9883), .Q(n10094), 
        .QN(n8223) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(n9024), .CK(CLK), .RN(n9883), .Q(n10095), 
        .QN(n8225) );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(n9016), .CK(CLK), .RN(n9883), .Q(n10103), 
        .QN(n8241) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(n9015), .CK(CLK), .RN(n9883), .Q(n10104), 
        .QN(n8243) );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(n9014), .CK(CLK), .RN(n9883), .Q(n10105), 
        .QN(n8245) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(n9012), .CK(CLK), .RN(n9883), .Q(n10011), 
        .QN(n2113) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(n9011), .CK(CLK), .RN(n9883), .Q(n10012), 
        .QN(n2121) );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(n9010), .CK(CLK), .RN(n9883), .Q(n10013), 
        .QN(n2129) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(n9009), .CK(CLK), .RN(n9883), .Q(n10014), 
        .QN(n2137) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(n9008), .CK(CLK), .RN(n9883), .Q(n10015), 
        .QN(n2145) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(n9007), .CK(CLK), .RN(n9883), .Q(n10016), 
        .QN(n2153) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(n9006), .CK(CLK), .RN(n9883), .Q(n10017), 
        .QN(n2161) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(n9005), .CK(CLK), .RN(n9883), .Q(n10018), 
        .QN(n2169) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(n9004), .CK(CLK), .RN(n9883), .Q(n10019), 
        .QN(n2177) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(n9003), .CK(CLK), .RN(n9883), .Q(n10020), 
        .QN(n2185) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(n9002), .CK(CLK), .RN(n9883), .Q(n10021), 
        .QN(n2193) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(n9001), .CK(CLK), .RN(n9883), .Q(n10022), 
        .QN(n2201) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(n9000), .CK(CLK), .RN(n9883), .Q(n10023), 
        .QN(n2209) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(n8999), .CK(CLK), .RN(n9883), .Q(n10024), 
        .QN(n2217) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(n8998), .CK(CLK), .RN(n9883), .Q(n10025), 
        .QN(n2225) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(n8997), .CK(CLK), .RN(n9883), .Q(n10026), 
        .QN(n2233) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(n8996), .CK(CLK), .RN(n9883), .Q(n10027), 
        .QN(n2241) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(n8995), .CK(CLK), .RN(n9883), .Q(n10028), 
        .QN(n2249) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(n8994), .CK(CLK), .RN(n9883), .Q(n10029), 
        .QN(n2257) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(n8993), .CK(CLK), .RN(n9883), .Q(n10030), 
        .QN(n2265) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(n8992), .CK(CLK), .RN(n9883), .Q(n10031), 
        .QN(n2273) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(n8984), .CK(CLK), .RN(n9883), .Q(n10039), 
        .QN(n2337) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(n8983), .CK(CLK), .RN(n9883), .Q(n10040), 
        .QN(n2345) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(n8982), .CK(CLK), .RN(n9883), .Q(n10041), 
        .QN(n2353) );
  DFFR_X1 \REGISTERS_reg[0][30]  ( .D(n8980), .CK(CLK), .RN(n9883), .Q(n9923), 
        .QN(n2112) );
  DFFR_X1 \REGISTERS_reg[0][29]  ( .D(n8979), .CK(CLK), .RN(n9883), .Q(n9924), 
        .QN(n2120) );
  DFFR_X1 \REGISTERS_reg[0][28]  ( .D(n8978), .CK(CLK), .RN(n9883), .Q(n9925), 
        .QN(n2128) );
  DFFR_X1 \REGISTERS_reg[0][27]  ( .D(n8977), .CK(CLK), .RN(n9883), .Q(n9926), 
        .QN(n2136) );
  DFFR_X1 \REGISTERS_reg[0][26]  ( .D(n8976), .CK(CLK), .RN(n9883), .Q(n9927), 
        .QN(n2144) );
  DFFR_X1 \REGISTERS_reg[0][25]  ( .D(n8975), .CK(CLK), .RN(n9883), .Q(n9928), 
        .QN(n2152) );
  DFFR_X1 \REGISTERS_reg[0][24]  ( .D(n8974), .CK(CLK), .RN(n9883), .Q(n9929), 
        .QN(n2160) );
  DFFR_X1 \REGISTERS_reg[0][23]  ( .D(n8973), .CK(CLK), .RN(n9883), .Q(n9930), 
        .QN(n2168) );
  DFFR_X1 \REGISTERS_reg[0][22]  ( .D(n8972), .CK(CLK), .RN(n9883), .Q(n9931), 
        .QN(n2176) );
  DFFR_X1 \REGISTERS_reg[0][21]  ( .D(n8971), .CK(CLK), .RN(n9883), .Q(n9932), 
        .QN(n2184) );
  DFFR_X1 \REGISTERS_reg[0][20]  ( .D(n8970), .CK(CLK), .RN(n9883), .Q(n9933), 
        .QN(n2192) );
  DFFR_X1 \REGISTERS_reg[0][19]  ( .D(n8969), .CK(CLK), .RN(n9883), .Q(n9934), 
        .QN(n2200) );
  DFFR_X1 \REGISTERS_reg[0][18]  ( .D(n8968), .CK(CLK), .RN(n9883), .Q(n9935), 
        .QN(n2208) );
  DFFR_X1 \REGISTERS_reg[0][17]  ( .D(n8967), .CK(CLK), .RN(n9883), .Q(n9936), 
        .QN(n2216) );
  DFFR_X1 \REGISTERS_reg[0][16]  ( .D(n8966), .CK(CLK), .RN(n9883), .Q(n9937), 
        .QN(n2224) );
  DFFR_X1 \REGISTERS_reg[0][15]  ( .D(n8965), .CK(CLK), .RN(n9883), .Q(n9938), 
        .QN(n2232) );
  DFFR_X1 \REGISTERS_reg[0][14]  ( .D(n8964), .CK(CLK), .RN(n9883), .Q(n9939), 
        .QN(n2240) );
  DFFR_X1 \REGISTERS_reg[0][13]  ( .D(n8963), .CK(CLK), .RN(n9883), .Q(n9940), 
        .QN(n2248) );
  DFFR_X1 \REGISTERS_reg[0][12]  ( .D(n8962), .CK(CLK), .RN(n9883), .Q(n9941), 
        .QN(n2256) );
  DFFR_X1 \REGISTERS_reg[0][11]  ( .D(n8961), .CK(CLK), .RN(n9883), .Q(n9942), 
        .QN(n2264) );
  DFFR_X1 \REGISTERS_reg[0][10]  ( .D(n8960), .CK(CLK), .RN(n9883), .Q(n9943), 
        .QN(n2272) );
  DFFR_X1 \REGISTERS_reg[0][2]  ( .D(n8952), .CK(CLK), .RN(n9883), .Q(n9951), 
        .QN(n2336) );
  DFFR_X1 \REGISTERS_reg[0][1]  ( .D(n8951), .CK(CLK), .RN(n9883), .Q(n9952), 
        .QN(n2344) );
  DFFR_X1 \REGISTERS_reg[0][0]  ( .D(n8950), .CK(CLK), .RN(n9883), .Q(n9953), 
        .QN(n2352) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(n3472), .CK(CLK), .RN(n9883), .Q(n10291), .QN(n8628) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(n3488), .CK(CLK), .RN(n9883), .Q(n10292), .QN(n8627) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(n3504), .CK(CLK), .RN(n9883), .Q(n10293), .QN(n8626) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(n3520), .CK(CLK), .RN(n9883), .Q(n10294), .QN(n8625) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(n3536), .CK(CLK), .RN(n9883), .Q(n10295), .QN(n8624) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(n3552), .CK(CLK), .RN(n9883), .Q(n10296), .QN(n8623) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(n3568), .CK(CLK), .RN(n9883), .Q(n10297), .QN(n8622) );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(n3584), .CK(CLK), .RN(n9883), .Q(n10298), .QN(n8621) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(n3600), .CK(CLK), .RN(n9883), .Q(n10299), .QN(n8620) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(n3616), .CK(CLK), .RN(n9883), .Q(n10300), .QN(n8619) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(n3632), .CK(CLK), .RN(n9883), .Q(n10301), .QN(n8618) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(n3648), .CK(CLK), .RN(n9883), .Q(n10302), .QN(n8617) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(n3664), .CK(CLK), .RN(n9883), .Q(n10303), .QN(n8616) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(n3680), .CK(CLK), .RN(n9883), .Q(n10304), .QN(n8615) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(n3696), .CK(CLK), .RN(n9883), .Q(n10305), .QN(n8614) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(n3712), .CK(CLK), .RN(n9883), .Q(n10306), .QN(n8613) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(n3728), .CK(CLK), .RN(n9883), .Q(n10307), .QN(n8612) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(n3744), .CK(CLK), .RN(n9883), .Q(n10308), .QN(n8611) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(n3760), .CK(CLK), .RN(n9883), .Q(n10309), .QN(n8610) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(n3776), .CK(CLK), .RN(n9883), .Q(n10310), .QN(n8609) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(n3792), .CK(CLK), .RN(n9883), .Q(n10311), .QN(n8608) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(n3920), .CK(CLK), .RN(n9883), .Q(n10319), 
        .QN(n8600) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(n3936), .CK(CLK), .RN(n9883), .Q(n10320), 
        .QN(n8599) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(n3952), .CK(CLK), .RN(n9883), .Q(n10321), 
        .QN(n8598) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(n3196), .CK(CLK), .RN(n9883), .QN(n8301) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(n3195), .CK(CLK), .RN(n9883), .QN(n8300) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(n3194), .CK(CLK), .RN(n9883), .QN(n8299) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(n3193), .CK(CLK), .RN(n9883), .QN(n8298) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(n3192), .CK(CLK), .RN(n9883), .QN(n8297) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(n3191), .CK(CLK), .RN(n9883), .QN(n8296) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(n3190), .CK(CLK), .RN(n9883), .QN(n8295) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(n3189), .CK(CLK), .RN(n9883), .QN(n8653) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(n3188), .CK(CLK), .RN(n9883), .QN(n8652) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(n3187), .CK(CLK), .RN(n9883), .QN(n8651) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(n3186), .CK(CLK), .RN(n9883), .QN(n8650) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(n3185), .CK(CLK), .RN(n9883), .QN(n8649) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(n3184), .CK(CLK), .RN(n9883), .QN(n8648) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(n3183), .CK(CLK), .RN(n9883), .QN(n8647) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(n3182), .CK(CLK), .RN(n9883), .QN(n8646) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(n3181), .CK(CLK), .RN(n9883), .QN(n8645) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(n3180), .CK(CLK), .RN(n9883), .QN(n8644) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(n3179), .CK(CLK), .RN(n9883), .QN(n8643) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(n3178), .CK(CLK), .RN(n9883), .QN(n8642) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(n3177), .CK(CLK), .RN(n9883), .QN(n8641) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(n3176), .CK(CLK), .RN(n9883), .QN(n8640) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(n3168), .CK(CLK), .RN(n9883), .QN(n8632)
         );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(n3167), .CK(CLK), .RN(n9883), .QN(n8631)
         );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(n3166), .CK(CLK), .RN(n9883), .QN(n8630)
         );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(n3228), .CK(CLK), .RN(n9883), .QN(n8684) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(n3227), .CK(CLK), .RN(n9883), .QN(n8683) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(n3226), .CK(CLK), .RN(n9883), .QN(n8682) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(n3225), .CK(CLK), .RN(n9883), .QN(n8681) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(n3224), .CK(CLK), .RN(n9883), .QN(n8680) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(n3223), .CK(CLK), .RN(n9883), .QN(n8679) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(n3222), .CK(CLK), .RN(n9883), .QN(n8678) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(n3221), .CK(CLK), .RN(n9883), .QN(n8677) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(n3220), .CK(CLK), .RN(n9883), .QN(n8676) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(n3219), .CK(CLK), .RN(n9883), .QN(n8675) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(n3218), .CK(CLK), .RN(n9883), .QN(n8674) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(n3217), .CK(CLK), .RN(n9883), .QN(n8673) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(n3216), .CK(CLK), .RN(n9883), .QN(n8672) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(n3215), .CK(CLK), .RN(n9883), .QN(n8671) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(n3214), .CK(CLK), .RN(n9883), .QN(n8670) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(n3213), .CK(CLK), .RN(n9883), .QN(n8669) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(n3212), .CK(CLK), .RN(n9883), .QN(n8668) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(n3211), .CK(CLK), .RN(n9883), .QN(n8667) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(n3210), .CK(CLK), .RN(n9883), .QN(n8666) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(n3209), .CK(CLK), .RN(n9883), .QN(n8665) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(n3208), .CK(CLK), .RN(n9883), .QN(n8664) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(n3200), .CK(CLK), .RN(n9883), .QN(n8656)
         );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(n3199), .CK(CLK), .RN(n9883), .QN(n8655)
         );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(n3198), .CK(CLK), .RN(n9883), .QN(n8654)
         );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(n3469), .CK(CLK), .RN(n9883), .Q(n10195), .QN(n8716) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(n3485), .CK(CLK), .RN(n9883), .Q(n10196), .QN(n8715) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(n3501), .CK(CLK), .RN(n9883), .Q(n10197), .QN(n8714) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(n3517), .CK(CLK), .RN(n9883), .Q(n10198), .QN(n8713) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(n3533), .CK(CLK), .RN(n9883), .Q(n10199), .QN(n8712) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(n3549), .CK(CLK), .RN(n9883), .Q(n10200), .QN(n8711) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(n3565), .CK(CLK), .RN(n9883), .Q(n10201), .QN(n8710) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(n3581), .CK(CLK), .RN(n9883), .Q(n10202), .QN(n8709) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(n3597), .CK(CLK), .RN(n9883), .Q(n10203), .QN(n8708) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(n3613), .CK(CLK), .RN(n9883), .Q(n10204), .QN(n8707) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(n3629), .CK(CLK), .RN(n9883), .Q(n10205), .QN(n8706) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(n3645), .CK(CLK), .RN(n9883), .Q(n10206), .QN(n8705) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(n3661), .CK(CLK), .RN(n9883), .Q(n10207), .QN(n8704) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(n3677), .CK(CLK), .RN(n9883), .Q(n10208), .QN(n8703) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(n3693), .CK(CLK), .RN(n9883), .Q(n10209), .QN(n8702) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(n3709), .CK(CLK), .RN(n9883), .Q(n10210), .QN(n8701) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(n3725), .CK(CLK), .RN(n9883), .Q(n10211), .QN(n8700) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(n3741), .CK(CLK), .RN(n9883), .Q(n10212), .QN(n8699) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(n3757), .CK(CLK), .RN(n9883), .Q(n10213), .QN(n8698) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(n3773), .CK(CLK), .RN(n9883), .Q(n10214), .QN(n8697) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(n3789), .CK(CLK), .RN(n9883), .Q(n10215), .QN(n8696) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(n3917), .CK(CLK), .RN(n9883), .Q(n10223), 
        .QN(n8688) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(n3933), .CK(CLK), .RN(n9883), .Q(n10224), 
        .QN(n8687) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(n3949), .CK(CLK), .RN(n9883), .Q(n10225), 
        .QN(n8686) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(n3260), .CK(CLK), .RN(n9883), .Q(n10579), .QN(n8293) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(n3259), .CK(CLK), .RN(n9883), .Q(n10580), .QN(n8292) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(n3258), .CK(CLK), .RN(n9883), .Q(n10581), .QN(n8291) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(n3257), .CK(CLK), .RN(n9883), .Q(n10582), .QN(n8290) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(n3256), .CK(CLK), .RN(n9883), .Q(n10583), .QN(n8289) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(n3255), .CK(CLK), .RN(n9883), .Q(n10584), .QN(n8288) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(n3254), .CK(CLK), .RN(n9883), .Q(n10585), .QN(n8287) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(n3253), .CK(CLK), .RN(n9883), .Q(n10170), .QN(n8741) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(n3252), .CK(CLK), .RN(n9883), .Q(n10171), .QN(n8740) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(n3251), .CK(CLK), .RN(n9883), .Q(n10172), .QN(n8739) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(n3250), .CK(CLK), .RN(n9883), .Q(n10173), .QN(n8738) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(n3249), .CK(CLK), .RN(n9883), .Q(n10174), .QN(n8737) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(n3248), .CK(CLK), .RN(n9883), .Q(n10175), .QN(n8736) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(n3247), .CK(CLK), .RN(n9883), .Q(n10176), .QN(n8735) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(n3246), .CK(CLK), .RN(n9883), .Q(n10177), .QN(n8734) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(n3245), .CK(CLK), .RN(n9883), .Q(n10178), .QN(n8733) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(n3244), .CK(CLK), .RN(n9883), .Q(n10179), .QN(n8732) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(n3243), .CK(CLK), .RN(n9883), .Q(n10180), .QN(n8731) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(n3242), .CK(CLK), .RN(n9883), .Q(n10181), .QN(n8730) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(n3241), .CK(CLK), .RN(n9883), .Q(n10182), .QN(n8729) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(n3240), .CK(CLK), .RN(n9883), .Q(n10183), .QN(n8728) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(n3232), .CK(CLK), .RN(n9883), .Q(n10191), 
        .QN(n8720) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(n3231), .CK(CLK), .RN(n9883), .Q(n10192), 
        .QN(n8719) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(n3230), .CK(CLK), .RN(n9883), .Q(n10193), 
        .QN(n8718) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(n3292), .CK(CLK), .RN(n9883), .Q(n10139), .QN(n8772) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(n3291), .CK(CLK), .RN(n9883), .Q(n10140), .QN(n8771) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(n3290), .CK(CLK), .RN(n9883), .Q(n10141), .QN(n8770) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(n3289), .CK(CLK), .RN(n9883), .Q(n10142), .QN(n8769) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(n3288), .CK(CLK), .RN(n9883), .Q(n10143), .QN(n8768) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(n3287), .CK(CLK), .RN(n9883), .Q(n10144), .QN(n8767) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(n3286), .CK(CLK), .RN(n9883), .Q(n10145), .QN(n8766) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(n3285), .CK(CLK), .RN(n9883), .Q(n10146), .QN(n8765) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(n3284), .CK(CLK), .RN(n9883), .Q(n10147), .QN(n8764) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(n3283), .CK(CLK), .RN(n9883), .Q(n10148), .QN(n8763) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(n3282), .CK(CLK), .RN(n9883), .Q(n10149), .QN(n8762) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(n3281), .CK(CLK), .RN(n9883), .Q(n10150), .QN(n8761) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(n3280), .CK(CLK), .RN(n9883), .Q(n10151), .QN(n8760) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(n3279), .CK(CLK), .RN(n9883), .Q(n10152), .QN(n8759) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(n3278), .CK(CLK), .RN(n9883), .Q(n10153), .QN(n8758) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(n3277), .CK(CLK), .RN(n9883), .Q(n10154), .QN(n8757) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(n3276), .CK(CLK), .RN(n9883), .Q(n10155), .QN(n8756) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(n3275), .CK(CLK), .RN(n9883), .Q(n10156), .QN(n8755) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(n3274), .CK(CLK), .RN(n9883), .Q(n10157), .QN(n8754) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(n3273), .CK(CLK), .RN(n9883), .Q(n10158), .QN(n8753) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(n3272), .CK(CLK), .RN(n9883), .Q(n10159), .QN(n8752) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(n3264), .CK(CLK), .RN(n9883), .Q(n10167), 
        .QN(n8744) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(n3263), .CK(CLK), .RN(n9883), .Q(n10168), 
        .QN(n8743) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(n3262), .CK(CLK), .RN(n9883), .Q(n10169), 
        .QN(n8742) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(n3468), .CK(CLK), .RN(n9883), .Q(n10107), 
        .QN(n2114) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(n3484), .CK(CLK), .RN(n9883), .Q(n10108), 
        .QN(n2122) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(n3500), .CK(CLK), .RN(n9883), .Q(n10109), 
        .QN(n2130) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(n3516), .CK(CLK), .RN(n9883), .Q(n10110), 
        .QN(n2138) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(n3532), .CK(CLK), .RN(n9883), .Q(n10111), 
        .QN(n2146) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(n3548), .CK(CLK), .RN(n9883), .Q(n10112), 
        .QN(n2154) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(n3564), .CK(CLK), .RN(n9883), .Q(n10113), 
        .QN(n2162) );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(n3580), .CK(CLK), .RN(n9883), .Q(n10114), 
        .QN(n2170) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(n3596), .CK(CLK), .RN(n9883), .Q(n10115), 
        .QN(n2178) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(n3612), .CK(CLK), .RN(n9883), .Q(n10116), 
        .QN(n2186) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(n3628), .CK(CLK), .RN(n9883), .Q(n10117), 
        .QN(n2194) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(n3644), .CK(CLK), .RN(n9883), .Q(n10118), 
        .QN(n2202) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(n3660), .CK(CLK), .RN(n9883), .Q(n10119), 
        .QN(n2210) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(n3676), .CK(CLK), .RN(n9883), .Q(n10120), 
        .QN(n2218) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(n3692), .CK(CLK), .RN(n9883), .Q(n10121), 
        .QN(n2226) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(n3708), .CK(CLK), .RN(n9883), .Q(n10122), 
        .QN(n2234) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(n3724), .CK(CLK), .RN(n9883), .Q(n10123), 
        .QN(n2242) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(n3740), .CK(CLK), .RN(n9883), .Q(n10124), 
        .QN(n2250) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(n3756), .CK(CLK), .RN(n9883), .Q(n10125), 
        .QN(n2258) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(n3772), .CK(CLK), .RN(n9883), .Q(n10126), 
        .QN(n2266) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(n3788), .CK(CLK), .RN(n9883), .Q(n10127), 
        .QN(n2274) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(n3916), .CK(CLK), .RN(n9883), .Q(n10135), 
        .QN(n2338) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(n3932), .CK(CLK), .RN(n9883), .Q(n10136), 
        .QN(n2346) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(n3948), .CK(CLK), .RN(n9883), .Q(n10137), 
        .QN(n2354) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(n3324), .CK(CLK), .RN(n9883), .QN(n8317)
         );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(n3323), .CK(CLK), .RN(n9883), .QN(n8316)
         );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(n3322), .CK(CLK), .RN(n9883), .QN(n8315)
         );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(n3321), .CK(CLK), .RN(n9883), .QN(n8314)
         );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(n3320), .CK(CLK), .RN(n9883), .QN(n8313)
         );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(n3319), .CK(CLK), .RN(n9883), .QN(n8312)
         );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(n3318), .CK(CLK), .RN(n9883), .QN(n8311)
         );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(n3317), .CK(CLK), .RN(n9883), .QN(n8797)
         );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(n3316), .CK(CLK), .RN(n9883), .QN(n8796)
         );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(n3315), .CK(CLK), .RN(n9883), .QN(n8795)
         );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(n3314), .CK(CLK), .RN(n9883), .QN(n8794)
         );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(n3313), .CK(CLK), .RN(n9883), .QN(n8793)
         );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(n3312), .CK(CLK), .RN(n9883), .QN(n8792)
         );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(n3311), .CK(CLK), .RN(n9883), .QN(n8791)
         );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(n3310), .CK(CLK), .RN(n9883), .QN(n8790)
         );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(n3309), .CK(CLK), .RN(n9883), .QN(n8789)
         );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(n3308), .CK(CLK), .RN(n9883), .QN(n8788)
         );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(n3307), .CK(CLK), .RN(n9883), .QN(n8787)
         );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(n3306), .CK(CLK), .RN(n9883), .QN(n8786)
         );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(n3305), .CK(CLK), .RN(n9883), .QN(n8785)
         );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(n3304), .CK(CLK), .RN(n9883), .QN(n8784)
         );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(n3296), .CK(CLK), .RN(n9883), .QN(n8776)
         );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(n3295), .CK(CLK), .RN(n9883), .QN(n8775)
         );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(n3294), .CK(CLK), .RN(n9883), .QN(n8774)
         );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(n3356), .CK(CLK), .RN(n9883), .QN(n8828)
         );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(n3355), .CK(CLK), .RN(n9883), .QN(n8827)
         );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(n3354), .CK(CLK), .RN(n9883), .QN(n8826)
         );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(n3353), .CK(CLK), .RN(n9883), .QN(n8825)
         );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(n3352), .CK(CLK), .RN(n9883), .QN(n8824)
         );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(n3351), .CK(CLK), .RN(n9883), .QN(n8823)
         );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(n3350), .CK(CLK), .RN(n9883), .QN(n8822)
         );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(n3349), .CK(CLK), .RN(n9883), .QN(n8821)
         );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(n3348), .CK(CLK), .RN(n9883), .QN(n8820)
         );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(n3347), .CK(CLK), .RN(n9883), .QN(n8819)
         );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(n3346), .CK(CLK), .RN(n9883), .QN(n8818)
         );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(n3345), .CK(CLK), .RN(n9883), .QN(n8817)
         );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(n3344), .CK(CLK), .RN(n9883), .QN(n8816)
         );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(n3343), .CK(CLK), .RN(n9883), .QN(n8815)
         );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(n3342), .CK(CLK), .RN(n9883), .QN(n8814)
         );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(n3341), .CK(CLK), .RN(n9883), .QN(n8813)
         );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(n3340), .CK(CLK), .RN(n9883), .QN(n8812)
         );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(n3339), .CK(CLK), .RN(n9883), .QN(n8811)
         );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(n3338), .CK(CLK), .RN(n9883), .QN(n8810)
         );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(n3337), .CK(CLK), .RN(n9883), .QN(n8809)
         );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(n3336), .CK(CLK), .RN(n9883), .QN(n8808)
         );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(n3328), .CK(CLK), .RN(n9883), .QN(n8800)
         );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(n3327), .CK(CLK), .RN(n9883), .QN(n8799)
         );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(n3326), .CK(CLK), .RN(n9883), .QN(n8798)
         );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(n3466), .CK(CLK), .RN(n9883), .Q(n10043), 
        .QN(n8860) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(n3482), .CK(CLK), .RN(n9883), .Q(n10044), 
        .QN(n8859) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(n3498), .CK(CLK), .RN(n9883), .Q(n10045), 
        .QN(n8858) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(n3514), .CK(CLK), .RN(n9883), .Q(n10046), 
        .QN(n8857) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(n3530), .CK(CLK), .RN(n9883), .Q(n10047), 
        .QN(n8856) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(n3546), .CK(CLK), .RN(n9883), .Q(n10048), 
        .QN(n8855) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(n3562), .CK(CLK), .RN(n9883), .Q(n10049), 
        .QN(n8854) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(n3578), .CK(CLK), .RN(n9883), .Q(n10050), 
        .QN(n8853) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(n3594), .CK(CLK), .RN(n9883), .Q(n10051), 
        .QN(n8852) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(n3610), .CK(CLK), .RN(n9883), .Q(n10052), 
        .QN(n8851) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(n3626), .CK(CLK), .RN(n9883), .Q(n10053), 
        .QN(n8850) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(n3642), .CK(CLK), .RN(n9883), .Q(n10054), 
        .QN(n8849) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(n3658), .CK(CLK), .RN(n9883), .Q(n10055), 
        .QN(n8848) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(n3674), .CK(CLK), .RN(n9883), .Q(n10056), 
        .QN(n8847) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(n3690), .CK(CLK), .RN(n9883), .Q(n10057), 
        .QN(n8846) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(n3706), .CK(CLK), .RN(n9883), .Q(n10058), 
        .QN(n8845) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(n3722), .CK(CLK), .RN(n9883), .Q(n10059), 
        .QN(n8844) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(n3738), .CK(CLK), .RN(n9883), .Q(n10060), 
        .QN(n8843) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(n3754), .CK(CLK), .RN(n9883), .Q(n10061), 
        .QN(n8842) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(n3770), .CK(CLK), .RN(n9883), .Q(n10062), 
        .QN(n8841) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(n3786), .CK(CLK), .RN(n9883), .Q(n10063), 
        .QN(n8840) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(n3914), .CK(CLK), .RN(n9883), .Q(n10071), 
        .QN(n8832) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(n3930), .CK(CLK), .RN(n9883), .Q(n10072), 
        .QN(n8831) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(n3946), .CK(CLK), .RN(n9883), .Q(n10073), 
        .QN(n8830) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(n3388), .CK(CLK), .RN(n9883), .Q(n10571), 
        .QN(n8309) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(n3387), .CK(CLK), .RN(n9883), .Q(n10572), 
        .QN(n8308) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(n3386), .CK(CLK), .RN(n9883), .Q(n10573), 
        .QN(n8307) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(n3385), .CK(CLK), .RN(n9883), .Q(n10574), 
        .QN(n8306) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(n3384), .CK(CLK), .RN(n9883), .Q(n10575), 
        .QN(n8305) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(n3383), .CK(CLK), .RN(n9883), .Q(n10576), 
        .QN(n8304) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(n3382), .CK(CLK), .RN(n9883), .Q(n10577), 
        .QN(n8303) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(n3381), .CK(CLK), .RN(n9883), .Q(n9986), 
        .QN(n8885) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(n3380), .CK(CLK), .RN(n9883), .Q(n9987), 
        .QN(n8884) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(n3379), .CK(CLK), .RN(n9883), .Q(n9988), 
        .QN(n8883) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(n3378), .CK(CLK), .RN(n9883), .Q(n9989), 
        .QN(n8882) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(n3377), .CK(CLK), .RN(n9883), .Q(n9990), 
        .QN(n8881) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(n3376), .CK(CLK), .RN(n9883), .Q(n9991), 
        .QN(n8880) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(n3375), .CK(CLK), .RN(n9883), .Q(n9992), 
        .QN(n8879) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(n3374), .CK(CLK), .RN(n9883), .Q(n9993), 
        .QN(n8878) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(n3373), .CK(CLK), .RN(n9883), .Q(n9994), 
        .QN(n8877) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(n3372), .CK(CLK), .RN(n9883), .Q(n9995), 
        .QN(n8876) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(n3371), .CK(CLK), .RN(n9883), .Q(n9996), 
        .QN(n8875) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(n3370), .CK(CLK), .RN(n9883), .Q(n9997), 
        .QN(n8874) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(n3369), .CK(CLK), .RN(n9883), .Q(n9998), 
        .QN(n8873) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(n3368), .CK(CLK), .RN(n9883), .Q(n9999), 
        .QN(n8872) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(n3360), .CK(CLK), .RN(n9883), .Q(n10007), 
        .QN(n8864) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(n3359), .CK(CLK), .RN(n9883), .Q(n10008), 
        .QN(n8863) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(n3358), .CK(CLK), .RN(n9883), .Q(n10009), 
        .QN(n8862) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(n3420), .CK(CLK), .RN(n9883), .QN(n8916)
         );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(n3419), .CK(CLK), .RN(n9883), .QN(n8915)
         );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(n3418), .CK(CLK), .RN(n9883), .QN(n8914)
         );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(n3417), .CK(CLK), .RN(n9883), .QN(n8913)
         );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(n3416), .CK(CLK), .RN(n9883), .QN(n8912)
         );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(n3415), .CK(CLK), .RN(n9883), .QN(n8911)
         );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(n3414), .CK(CLK), .RN(n9883), .QN(n8910)
         );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(n3413), .CK(CLK), .RN(n9883), .QN(n8909)
         );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(n3412), .CK(CLK), .RN(n9883), .QN(n8908)
         );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(n3411), .CK(CLK), .RN(n9883), .QN(n8907)
         );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(n3410), .CK(CLK), .RN(n9883), .QN(n8906)
         );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(n3409), .CK(CLK), .RN(n9883), .QN(n8905)
         );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(n3408), .CK(CLK), .RN(n9883), .QN(n8904)
         );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(n3407), .CK(CLK), .RN(n9883), .QN(n8903)
         );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(n3406), .CK(CLK), .RN(n9883), .QN(n8902)
         );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(n3405), .CK(CLK), .RN(n9883), .QN(n8901)
         );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(n3404), .CK(CLK), .RN(n9883), .QN(n8900)
         );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(n3403), .CK(CLK), .RN(n9883), .QN(n8899)
         );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(n3402), .CK(CLK), .RN(n9883), .QN(n8898)
         );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(n3401), .CK(CLK), .RN(n9883), .QN(n8897)
         );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(n3400), .CK(CLK), .RN(n9883), .QN(n8896)
         );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(n3392), .CK(CLK), .RN(n9883), .QN(n8888)
         );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(n3391), .CK(CLK), .RN(n9883), .QN(n8887)
         );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(n3390), .CK(CLK), .RN(n9883), .QN(n8886)
         );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(n3464), .CK(CLK), .RN(n9883), .Q(n9955), 
        .QN(n8948) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(n3480), .CK(CLK), .RN(n9883), .Q(n9956), 
        .QN(n8947) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(n3496), .CK(CLK), .RN(n9883), .Q(n9957), 
        .QN(n8946) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(n3512), .CK(CLK), .RN(n9883), .Q(n9958), 
        .QN(n8945) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(n3528), .CK(CLK), .RN(n9883), .Q(n9959), 
        .QN(n8944) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(n3544), .CK(CLK), .RN(n9883), .Q(n9960), 
        .QN(n8943) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(n3560), .CK(CLK), .RN(n9883), .Q(n9961), 
        .QN(n8942) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(n3576), .CK(CLK), .RN(n9883), .Q(n9962), 
        .QN(n8941) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(n3592), .CK(CLK), .RN(n9883), .Q(n9963), 
        .QN(n8940) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(n3608), .CK(CLK), .RN(n9883), .Q(n9964), 
        .QN(n8939) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(n3624), .CK(CLK), .RN(n9883), .Q(n9965), 
        .QN(n8938) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(n3640), .CK(CLK), .RN(n9883), .Q(n9966), 
        .QN(n8937) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(n3656), .CK(CLK), .RN(n9883), .Q(n9967), 
        .QN(n8936) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(n3672), .CK(CLK), .RN(n9883), .Q(n9968), 
        .QN(n8935) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(n3688), .CK(CLK), .RN(n9883), .Q(n9969), 
        .QN(n8934) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(n3704), .CK(CLK), .RN(n9883), .Q(n9970), 
        .QN(n8933) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(n3720), .CK(CLK), .RN(n9883), .Q(n9971), 
        .QN(n8932) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(n3736), .CK(CLK), .RN(n9883), .Q(n9972), 
        .QN(n8931) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(n3752), .CK(CLK), .RN(n9883), .Q(n9973), 
        .QN(n8930) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(n3768), .CK(CLK), .RN(n9883), .Q(n9974), 
        .QN(n8929) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(n3784), .CK(CLK), .RN(n9883), .Q(n9975), 
        .QN(n8928) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(n3912), .CK(CLK), .RN(n9883), .Q(n9983), 
        .QN(n8920) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(n3928), .CK(CLK), .RN(n9883), .Q(n9984), 
        .QN(n8919) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(n3944), .CK(CLK), .RN(n9883), .Q(n9985), 
        .QN(n8918) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(n9204), .CK(CLK), .RN(n9878), .Q(n10347), .QN(n2109) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(n9203), .CK(CLK), .RN(n9878), .Q(n10348), .QN(n2117) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(n9202), .CK(CLK), .RN(n9878), .Q(n10349), .QN(n2125) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(n9201), .CK(CLK), .RN(n9878), .Q(n10350), .QN(n2133) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(n9200), .CK(CLK), .RN(n9883), .Q(n10351), .QN(n2141) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(n9199), .CK(CLK), .RN(n9878), .Q(n10352), .QN(n2149) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(n9198), .CK(CLK), .RN(n9878), .Q(n10353), .QN(n2157) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(n9183), .CK(CLK), .RN(n9883), .Q(n10368), 
        .QN(n2277) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(n9197), .CK(CLK), .RN(n9877), .Q(n10354), .QN(n2165) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(n9196), .CK(CLK), .RN(n9877), .Q(n10355), .QN(n2173) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(n9195), .CK(CLK), .RN(n9877), .Q(n10356), .QN(n2181) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(n9194), .CK(CLK), .RN(n9877), .Q(n10357), .QN(n2189) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(n9193), .CK(CLK), .RN(n9883), .Q(n10358), .QN(n2197) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(n9192), .CK(CLK), .RN(n9883), .Q(n10359), .QN(n2205) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(n9191), .CK(CLK), .RN(n9883), .Q(n10360), .QN(n2213) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(n9190), .CK(CLK), .RN(n9877), .Q(n10361), .QN(n2221) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(n9189), .CK(CLK), .RN(n9877), .Q(n10362), .QN(n2229) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(n9188), .CK(CLK), .RN(n9883), .Q(n10363), .QN(n2237) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(n9187), .CK(CLK), .RN(n9883), .Q(n10364), .QN(n2245) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(n9186), .CK(CLK), .RN(n9883), .Q(n10365), .QN(n2253) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(n9185), .CK(CLK), .RN(n9882), .Q(n10366), .QN(n2261) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(n9184), .CK(CLK), .RN(n9883), .Q(n10367), .QN(n2269) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(n9182), .CK(CLK), .RN(n9883), .Q(n10369), 
        .QN(n2285) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(n9181), .CK(CLK), .RN(n9883), .Q(n10370), 
        .QN(n2293) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(n9180), .CK(CLK), .RN(n9883), .Q(n10371), 
        .QN(n2301) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(n9179), .CK(CLK), .RN(n9883), .Q(n10372), 
        .QN(n2309) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(n9178), .CK(CLK), .RN(n9883), .Q(n10373), 
        .QN(n2317) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(n9177), .CK(CLK), .RN(n9877), .Q(n10374), 
        .QN(n2325) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(n9176), .CK(CLK), .RN(n9883), .Q(n10375), 
        .QN(n2333) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(n9175), .CK(CLK), .RN(n9883), .Q(n10376), 
        .QN(n2341) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(n9174), .CK(CLK), .RN(n9877), .Q(n10377), 
        .QN(n2349) );
  AND2_X1 U2 ( .A1(n822), .A2(n816), .ZN(n9207) );
  AND2_X1 U3 ( .A1(n819), .A2(n816), .ZN(n9208) );
  AND2_X1 U4 ( .A1(n824), .A2(n821), .ZN(n9209) );
  AND2_X1 U5 ( .A1(n827), .A2(n816), .ZN(n9210) );
  AND2_X1 U6 ( .A1(n824), .A2(n816), .ZN(n9211) );
  AND2_X1 U7 ( .A1(n827), .A2(n821), .ZN(n9212) );
  AND2_X1 U8 ( .A1(n847), .A2(n826), .ZN(n9213) );
  AND2_X1 U9 ( .A1(n842), .A2(n816), .ZN(n9214) );
  AND2_X1 U10 ( .A1(n842), .A2(n830), .ZN(n9215) );
  AND2_X1 U11 ( .A1(n847), .A2(n816), .ZN(n9216) );
  AND2_X1 U12 ( .A1(n847), .A2(n830), .ZN(n9217) );
  AND2_X1 U13 ( .A1(n842), .A2(n821), .ZN(n9218) );
  AND2_X1 U14 ( .A1(n845), .A2(n816), .ZN(n9219) );
  AND2_X1 U15 ( .A1(n845), .A2(n826), .ZN(n9220) );
  AND2_X1 U16 ( .A1(n845), .A2(n830), .ZN(n9221) );
  AND2_X1 U17 ( .A1(n847), .A2(n821), .ZN(n9222) );
  AND2_X1 U18 ( .A1(n845), .A2(n821), .ZN(n9223) );
  AND2_X1 U19 ( .A1(n842), .A2(n826), .ZN(n9224) );
  AND2_X1 U20 ( .A1(n821), .A2(n819), .ZN(n9225) );
  AND2_X1 U21 ( .A1(n826), .A2(n822), .ZN(n9226) );
  AND2_X1 U22 ( .A1(n830), .A2(n827), .ZN(n9227) );
  AND2_X1 U23 ( .A1(n821), .A2(n817), .ZN(n9228) );
  AND2_X1 U24 ( .A1(n830), .A2(n824), .ZN(n9229) );
  AND2_X1 U25 ( .A1(n830), .A2(n822), .ZN(n9230) );
  AND2_X1 U26 ( .A1(n821), .A2(n822), .ZN(n9231) );
  AND2_X1 U27 ( .A1(n826), .A2(n819), .ZN(n9232) );
  AND2_X1 U28 ( .A1(n826), .A2(n824), .ZN(n9233) );
  AND2_X1 U29 ( .A1(n826), .A2(n827), .ZN(n9234) );
  AND2_X1 U30 ( .A1(n826), .A2(n817), .ZN(n9235) );
  AND2_X1 U31 ( .A1(n830), .A2(n817), .ZN(n9236) );
  AND2_X1 U32 ( .A1(n830), .A2(n819), .ZN(n9237) );
  INV_X32 U33 ( .A(n9876), .ZN(n9883) );
  CLKBUF_X1 U34 ( .A(RESET), .Z(n9876) );
  INV_X1 U35 ( .A(n9646), .ZN(n9636) );
  INV_X1 U36 ( .A(n9646), .ZN(n9637) );
  INV_X1 U37 ( .A(n9558), .ZN(n9549) );
  INV_X1 U38 ( .A(n9536), .ZN(n9526) );
  INV_X1 U39 ( .A(n9536), .ZN(n9527) );
  INV_X1 U40 ( .A(n9855), .ZN(n9846) );
  INV_X1 U41 ( .A(n9547), .ZN(n9537) );
  INV_X1 U42 ( .A(n9547), .ZN(n9538) );
  INV_X1 U43 ( .A(n9855), .ZN(n9845) );
  INV_X1 U44 ( .A(n9844), .ZN(n9835) );
  INV_X1 U45 ( .A(n9844), .ZN(n9834) );
  INV_X1 U46 ( .A(n9789), .ZN(n9780) );
  INV_X1 U47 ( .A(n9789), .ZN(n9779) );
  INV_X1 U48 ( .A(n9778), .ZN(n9769) );
  INV_X1 U49 ( .A(n9778), .ZN(n9768) );
  INV_X1 U50 ( .A(n9767), .ZN(n9758) );
  INV_X1 U51 ( .A(n9767), .ZN(n9757) );
  INV_X1 U52 ( .A(n9756), .ZN(n9747) );
  INV_X1 U53 ( .A(n9756), .ZN(n9746) );
  INV_X1 U54 ( .A(n9558), .ZN(n9548) );
  INV_X1 U55 ( .A(n9569), .ZN(n9559) );
  INV_X1 U56 ( .A(n9569), .ZN(n9560) );
  INV_X1 U57 ( .A(n9745), .ZN(n9736) );
  INV_X1 U58 ( .A(n9745), .ZN(n9735) );
  INV_X1 U59 ( .A(n9580), .ZN(n9570) );
  INV_X1 U60 ( .A(n9580), .ZN(n9571) );
  INV_X1 U61 ( .A(n9591), .ZN(n9581) );
  INV_X1 U62 ( .A(n9591), .ZN(n9582) );
  INV_X1 U63 ( .A(n9734), .ZN(n9725) );
  INV_X1 U64 ( .A(n9734), .ZN(n9724) );
  INV_X1 U65 ( .A(n9866), .ZN(n9856) );
  INV_X1 U66 ( .A(n9866), .ZN(n9857) );
  INV_X1 U67 ( .A(n9602), .ZN(n9592) );
  INV_X1 U68 ( .A(n9602), .ZN(n9593) );
  INV_X1 U69 ( .A(n9613), .ZN(n9603) );
  INV_X1 U70 ( .A(n9613), .ZN(n9604) );
  INV_X1 U71 ( .A(n9833), .ZN(n9823) );
  INV_X1 U72 ( .A(n9833), .ZN(n9824) );
  INV_X1 U73 ( .A(n9723), .ZN(n9714) );
  INV_X1 U74 ( .A(n9723), .ZN(n9713) );
  INV_X1 U75 ( .A(n9624), .ZN(n9614) );
  INV_X1 U76 ( .A(n9624), .ZN(n9615) );
  INV_X1 U77 ( .A(n9635), .ZN(n9625) );
  INV_X1 U78 ( .A(n9635), .ZN(n9626) );
  INV_X1 U79 ( .A(n9712), .ZN(n9703) );
  INV_X1 U80 ( .A(n9712), .ZN(n9702) );
  INV_X1 U81 ( .A(n9822), .ZN(n9812) );
  INV_X1 U82 ( .A(n9822), .ZN(n9813) );
  INV_X1 U83 ( .A(n9657), .ZN(n9647) );
  INV_X1 U84 ( .A(n9657), .ZN(n9648) );
  INV_X1 U85 ( .A(n9701), .ZN(n9692) );
  INV_X1 U86 ( .A(n9701), .ZN(n9691) );
  INV_X1 U87 ( .A(n9811), .ZN(n9801) );
  INV_X1 U88 ( .A(n9811), .ZN(n9802) );
  INV_X1 U89 ( .A(n9668), .ZN(n9658) );
  INV_X1 U90 ( .A(n9668), .ZN(n9659) );
  INV_X1 U91 ( .A(n9679), .ZN(n9669) );
  INV_X1 U92 ( .A(n9679), .ZN(n9670) );
  INV_X1 U93 ( .A(n9690), .ZN(n9681) );
  INV_X1 U94 ( .A(n9690), .ZN(n9680) );
  INV_X1 U95 ( .A(n9800), .ZN(n9790) );
  INV_X1 U96 ( .A(n9800), .ZN(n9791) );
  BUF_X1 U97 ( .A(n9229), .Z(n9646) );
  BUF_X1 U98 ( .A(n9229), .Z(n9639) );
  BUF_X1 U99 ( .A(n9229), .Z(n9638) );
  BUF_X1 U100 ( .A(n9643), .Z(n9645) );
  BUF_X1 U101 ( .A(n9642), .Z(n9644) );
  BUF_X1 U102 ( .A(n9229), .Z(n9643) );
  BUF_X1 U103 ( .A(n9229), .Z(n9642) );
  BUF_X1 U104 ( .A(n9229), .Z(n9641) );
  BUF_X1 U105 ( .A(n9229), .Z(n9640) );
  INV_X1 U106 ( .A(n9875), .ZN(n9867) );
  INV_X1 U107 ( .A(n9875), .ZN(n9868) );
  BUF_X1 U108 ( .A(n9210), .Z(n9745) );
  BUF_X1 U109 ( .A(n9207), .Z(n9591) );
  BUF_X1 U110 ( .A(n9208), .Z(n9866) );
  BUF_X1 U111 ( .A(n9222), .Z(n9536) );
  BUF_X1 U112 ( .A(n9223), .Z(n9547) );
  BUF_X1 U113 ( .A(n9209), .Z(n9844) );
  BUF_X1 U114 ( .A(n9212), .Z(n9789) );
  BUF_X1 U115 ( .A(n9218), .Z(n9767) );
  BUF_X1 U116 ( .A(n9211), .Z(n9558) );
  BUF_X1 U117 ( .A(n9216), .Z(n9569) );
  BUF_X1 U118 ( .A(n9219), .Z(n9580) );
  BUF_X1 U119 ( .A(n9214), .Z(n9734) );
  BUF_X1 U120 ( .A(n9213), .Z(n9613) );
  BUF_X1 U121 ( .A(n9220), .Z(n9624) );
  BUF_X1 U122 ( .A(n9224), .Z(n9712) );
  BUF_X1 U123 ( .A(n9217), .Z(n9657) );
  BUF_X1 U124 ( .A(n9221), .Z(n9668) );
  BUF_X1 U125 ( .A(n9215), .Z(n9690) );
  BUF_X1 U126 ( .A(n9231), .Z(n9855) );
  BUF_X1 U127 ( .A(n9228), .Z(n9778) );
  BUF_X1 U128 ( .A(n9225), .Z(n9756) );
  BUF_X1 U129 ( .A(n9233), .Z(n9602) );
  BUF_X1 U130 ( .A(n9234), .Z(n9833) );
  BUF_X1 U131 ( .A(n9235), .Z(n9723) );
  BUF_X1 U132 ( .A(n9226), .Z(n9635) );
  BUF_X1 U133 ( .A(n9232), .Z(n9822) );
  BUF_X1 U134 ( .A(n9227), .Z(n9701) );
  BUF_X1 U135 ( .A(n9236), .Z(n9811) );
  BUF_X1 U136 ( .A(n9230), .Z(n9679) );
  BUF_X1 U137 ( .A(n9237), .Z(n9800) );
  BUF_X1 U138 ( .A(n9211), .Z(n9555) );
  BUF_X1 U139 ( .A(n9211), .Z(n9554) );
  BUF_X1 U140 ( .A(n9211), .Z(n9553) );
  BUF_X1 U141 ( .A(n9211), .Z(n9552) );
  BUF_X1 U142 ( .A(n9209), .Z(n9838) );
  BUF_X1 U143 ( .A(n9209), .Z(n9840) );
  BUF_X1 U144 ( .A(n9840), .Z(n9842) );
  BUF_X1 U145 ( .A(n9839), .Z(n9843) );
  BUF_X1 U146 ( .A(n9212), .Z(n9783) );
  BUF_X1 U147 ( .A(n9212), .Z(n9784) );
  BUF_X1 U148 ( .A(n9212), .Z(n9785) );
  BUF_X1 U149 ( .A(n9212), .Z(n9786) );
  BUF_X1 U150 ( .A(n9784), .Z(n9787) );
  BUF_X1 U151 ( .A(n9785), .Z(n9788) );
  BUF_X1 U152 ( .A(n9210), .Z(n9742) );
  BUF_X1 U153 ( .A(n9585), .Z(n9589) );
  BUF_X1 U154 ( .A(n9207), .Z(n9588) );
  BUF_X1 U155 ( .A(n9207), .Z(n9587) );
  BUF_X1 U156 ( .A(n9207), .Z(n9586) );
  BUF_X1 U157 ( .A(n9207), .Z(n9585) );
  BUF_X1 U158 ( .A(n9207), .Z(n9584) );
  BUF_X1 U159 ( .A(n9207), .Z(n9583) );
  BUF_X1 U160 ( .A(n9860), .Z(n9865) );
  BUF_X1 U161 ( .A(n9859), .Z(n9864) );
  BUF_X1 U162 ( .A(n9208), .Z(n9863) );
  BUF_X1 U163 ( .A(n9208), .Z(n9862) );
  BUF_X1 U164 ( .A(n9208), .Z(n9861) );
  BUF_X1 U165 ( .A(n9208), .Z(n9860) );
  BUF_X1 U166 ( .A(n9208), .Z(n9859) );
  BUF_X1 U167 ( .A(n9208), .Z(n9858) );
  BUF_X1 U168 ( .A(n9530), .Z(n9535) );
  BUF_X1 U169 ( .A(n9533), .Z(n9534) );
  BUF_X1 U170 ( .A(n9222), .Z(n9533) );
  BUF_X1 U171 ( .A(n9222), .Z(n9532) );
  BUF_X1 U172 ( .A(n9222), .Z(n9531) );
  BUF_X1 U173 ( .A(n9222), .Z(n9530) );
  BUF_X1 U174 ( .A(n9541), .Z(n9546) );
  BUF_X1 U175 ( .A(n9544), .Z(n9545) );
  BUF_X1 U176 ( .A(n9223), .Z(n9544) );
  BUF_X1 U177 ( .A(n9223), .Z(n9543) );
  BUF_X1 U178 ( .A(n9223), .Z(n9542) );
  BUF_X1 U179 ( .A(n9223), .Z(n9541) );
  BUF_X1 U180 ( .A(n9220), .Z(n9617) );
  BUF_X1 U181 ( .A(n9220), .Z(n9616) );
  BUF_X1 U182 ( .A(n9221), .Z(n9661) );
  BUF_X1 U183 ( .A(n9221), .Z(n9660) );
  BUF_X1 U184 ( .A(n9219), .Z(n9573) );
  BUF_X1 U185 ( .A(n9219), .Z(n9572) );
  BUF_X1 U186 ( .A(n9211), .Z(n9551) );
  BUF_X1 U187 ( .A(n9211), .Z(n9550) );
  BUF_X1 U188 ( .A(n9222), .Z(n9529) );
  BUF_X1 U189 ( .A(n9222), .Z(n9528) );
  BUF_X1 U190 ( .A(n9223), .Z(n9540) );
  BUF_X1 U191 ( .A(n9223), .Z(n9539) );
  BUF_X1 U192 ( .A(n9209), .Z(n9836) );
  BUF_X1 U193 ( .A(n9209), .Z(n9837) );
  BUF_X1 U194 ( .A(n9209), .Z(n9839) );
  BUF_X1 U195 ( .A(n9209), .Z(n9841) );
  BUF_X1 U196 ( .A(n9212), .Z(n9781) );
  BUF_X1 U197 ( .A(n9212), .Z(n9782) );
  BUF_X1 U198 ( .A(n9218), .Z(n9759) );
  BUF_X1 U199 ( .A(n9218), .Z(n9760) );
  BUF_X1 U200 ( .A(n9218), .Z(n9761) );
  BUF_X1 U201 ( .A(n9218), .Z(n9762) );
  BUF_X1 U202 ( .A(n9218), .Z(n9763) );
  BUF_X1 U203 ( .A(n9218), .Z(n9764) );
  BUF_X1 U204 ( .A(n9762), .Z(n9765) );
  BUF_X1 U205 ( .A(n9763), .Z(n9766) );
  BUF_X1 U206 ( .A(n9552), .Z(n9557) );
  BUF_X1 U207 ( .A(n9555), .Z(n9556) );
  BUF_X1 U208 ( .A(n9563), .Z(n9568) );
  BUF_X1 U209 ( .A(n9566), .Z(n9567) );
  BUF_X1 U210 ( .A(n9216), .Z(n9566) );
  BUF_X1 U211 ( .A(n9216), .Z(n9565) );
  BUF_X1 U212 ( .A(n9216), .Z(n9564) );
  BUF_X1 U213 ( .A(n9216), .Z(n9563) );
  BUF_X1 U214 ( .A(n9216), .Z(n9562) );
  BUF_X1 U215 ( .A(n9216), .Z(n9561) );
  BUF_X1 U216 ( .A(n9210), .Z(n9737) );
  BUF_X1 U217 ( .A(n9210), .Z(n9738) );
  BUF_X1 U218 ( .A(n9210), .Z(n9739) );
  BUF_X1 U219 ( .A(n9210), .Z(n9740) );
  BUF_X1 U220 ( .A(n9210), .Z(n9741) );
  BUF_X1 U221 ( .A(n9742), .Z(n9743) );
  BUF_X1 U222 ( .A(n9740), .Z(n9744) );
  BUF_X1 U223 ( .A(n9588), .Z(n9590) );
  BUF_X1 U224 ( .A(n9574), .Z(n9579) );
  BUF_X1 U225 ( .A(n9577), .Z(n9578) );
  BUF_X1 U226 ( .A(n9219), .Z(n9577) );
  BUF_X1 U227 ( .A(n9219), .Z(n9576) );
  BUF_X1 U228 ( .A(n9219), .Z(n9575) );
  BUF_X1 U229 ( .A(n9219), .Z(n9574) );
  BUF_X1 U230 ( .A(n9214), .Z(n9726) );
  BUF_X1 U231 ( .A(n9214), .Z(n9727) );
  BUF_X1 U232 ( .A(n9214), .Z(n9728) );
  BUF_X1 U233 ( .A(n9214), .Z(n9729) );
  BUF_X1 U234 ( .A(n9214), .Z(n9730) );
  BUF_X1 U235 ( .A(n9214), .Z(n9731) );
  BUF_X1 U236 ( .A(n9726), .Z(n9732) );
  BUF_X1 U237 ( .A(n9727), .Z(n9733) );
  BUF_X1 U238 ( .A(n9610), .Z(n9612) );
  BUF_X1 U239 ( .A(n9609), .Z(n9611) );
  BUF_X1 U240 ( .A(n9213), .Z(n9610) );
  BUF_X1 U241 ( .A(n9213), .Z(n9609) );
  BUF_X1 U242 ( .A(n9213), .Z(n9608) );
  BUF_X1 U243 ( .A(n9213), .Z(n9607) );
  BUF_X1 U244 ( .A(n9213), .Z(n9606) );
  BUF_X1 U245 ( .A(n9213), .Z(n9605) );
  BUF_X1 U246 ( .A(n9617), .Z(n9623) );
  BUF_X1 U247 ( .A(n9616), .Z(n9622) );
  BUF_X1 U248 ( .A(n9220), .Z(n9621) );
  BUF_X1 U249 ( .A(n9220), .Z(n9620) );
  BUF_X1 U250 ( .A(n9220), .Z(n9619) );
  BUF_X1 U251 ( .A(n9220), .Z(n9618) );
  BUF_X1 U252 ( .A(n9224), .Z(n9704) );
  BUF_X1 U253 ( .A(n9224), .Z(n9705) );
  BUF_X1 U254 ( .A(n9224), .Z(n9706) );
  BUF_X1 U255 ( .A(n9224), .Z(n9707) );
  BUF_X1 U256 ( .A(n9224), .Z(n9708) );
  BUF_X1 U257 ( .A(n9224), .Z(n9709) );
  BUF_X1 U258 ( .A(n9707), .Z(n9710) );
  BUF_X1 U259 ( .A(n9708), .Z(n9711) );
  BUF_X1 U260 ( .A(n9651), .Z(n9656) );
  BUF_X1 U261 ( .A(n9650), .Z(n9655) );
  BUF_X1 U262 ( .A(n9217), .Z(n9654) );
  BUF_X1 U263 ( .A(n9217), .Z(n9653) );
  BUF_X1 U264 ( .A(n9217), .Z(n9652) );
  BUF_X1 U265 ( .A(n9217), .Z(n9651) );
  BUF_X1 U266 ( .A(n9217), .Z(n9650) );
  BUF_X1 U267 ( .A(n9217), .Z(n9649) );
  BUF_X1 U268 ( .A(n9661), .Z(n9667) );
  BUF_X1 U269 ( .A(n9660), .Z(n9666) );
  BUF_X1 U270 ( .A(n9221), .Z(n9665) );
  BUF_X1 U271 ( .A(n9221), .Z(n9664) );
  BUF_X1 U272 ( .A(n9221), .Z(n9663) );
  BUF_X1 U273 ( .A(n9221), .Z(n9662) );
  BUF_X1 U274 ( .A(n9215), .Z(n9682) );
  BUF_X1 U275 ( .A(n9215), .Z(n9683) );
  BUF_X1 U276 ( .A(n9215), .Z(n9684) );
  BUF_X1 U277 ( .A(n9215), .Z(n9685) );
  BUF_X1 U278 ( .A(n9215), .Z(n9686) );
  BUF_X1 U279 ( .A(n9215), .Z(n9687) );
  BUF_X1 U280 ( .A(n9685), .Z(n9688) );
  BUF_X1 U281 ( .A(n9686), .Z(n9689) );
  BUF_X1 U282 ( .A(n9231), .Z(n9847) );
  BUF_X1 U283 ( .A(n9231), .Z(n9848) );
  BUF_X1 U284 ( .A(n9231), .Z(n9849) );
  BUF_X1 U285 ( .A(n9231), .Z(n9850) );
  BUF_X1 U286 ( .A(n9231), .Z(n9851) );
  BUF_X1 U287 ( .A(n9231), .Z(n9852) );
  BUF_X1 U288 ( .A(n9233), .Z(n9595) );
  BUF_X1 U289 ( .A(n9233), .Z(n9594) );
  BUF_X1 U290 ( .A(n9850), .Z(n9853) );
  BUF_X1 U291 ( .A(n9851), .Z(n9854) );
  BUF_X1 U292 ( .A(n9228), .Z(n9770) );
  BUF_X1 U293 ( .A(n9228), .Z(n9771) );
  BUF_X1 U294 ( .A(n9228), .Z(n9772) );
  BUF_X1 U295 ( .A(n9228), .Z(n9773) );
  BUF_X1 U296 ( .A(n9228), .Z(n9774) );
  BUF_X1 U297 ( .A(n9228), .Z(n9775) );
  BUF_X1 U298 ( .A(n9773), .Z(n9776) );
  BUF_X1 U299 ( .A(n9774), .Z(n9777) );
  BUF_X1 U300 ( .A(n9225), .Z(n9748) );
  BUF_X1 U301 ( .A(n9225), .Z(n9749) );
  BUF_X1 U302 ( .A(n9225), .Z(n9750) );
  BUF_X1 U303 ( .A(n9225), .Z(n9751) );
  BUF_X1 U304 ( .A(n9225), .Z(n9752) );
  BUF_X1 U305 ( .A(n9225), .Z(n9753) );
  BUF_X1 U306 ( .A(n9751), .Z(n9754) );
  BUF_X1 U307 ( .A(n9752), .Z(n9755) );
  BUF_X1 U308 ( .A(n9599), .Z(n9601) );
  BUF_X1 U309 ( .A(n9598), .Z(n9600) );
  BUF_X1 U310 ( .A(n9233), .Z(n9599) );
  BUF_X1 U311 ( .A(n9233), .Z(n9598) );
  BUF_X1 U312 ( .A(n9233), .Z(n9597) );
  BUF_X1 U313 ( .A(n9233), .Z(n9596) );
  BUF_X1 U314 ( .A(n9827), .Z(n9832) );
  BUF_X1 U315 ( .A(n9826), .Z(n9831) );
  BUF_X1 U316 ( .A(n9234), .Z(n9830) );
  BUF_X1 U317 ( .A(n9234), .Z(n9829) );
  BUF_X1 U318 ( .A(n9234), .Z(n9828) );
  BUF_X1 U319 ( .A(n9234), .Z(n9827) );
  BUF_X1 U320 ( .A(n9234), .Z(n9826) );
  BUF_X1 U321 ( .A(n9234), .Z(n9825) );
  BUF_X1 U322 ( .A(n9235), .Z(n9715) );
  BUF_X1 U323 ( .A(n9235), .Z(n9716) );
  BUF_X1 U324 ( .A(n9235), .Z(n9717) );
  BUF_X1 U325 ( .A(n9235), .Z(n9718) );
  BUF_X1 U326 ( .A(n9235), .Z(n9719) );
  BUF_X1 U327 ( .A(n9235), .Z(n9720) );
  BUF_X1 U328 ( .A(n9718), .Z(n9721) );
  BUF_X1 U329 ( .A(n9719), .Z(n9722) );
  BUF_X1 U330 ( .A(n9629), .Z(n9634) );
  BUF_X1 U331 ( .A(n9628), .Z(n9633) );
  BUF_X1 U332 ( .A(n9226), .Z(n9632) );
  BUF_X1 U333 ( .A(n9226), .Z(n9631) );
  BUF_X1 U334 ( .A(n9226), .Z(n9630) );
  BUF_X1 U335 ( .A(n9226), .Z(n9629) );
  BUF_X1 U336 ( .A(n9226), .Z(n9628) );
  BUF_X1 U337 ( .A(n9226), .Z(n9627) );
  BUF_X1 U338 ( .A(n9819), .Z(n9821) );
  BUF_X1 U339 ( .A(n9818), .Z(n9820) );
  BUF_X1 U340 ( .A(n9232), .Z(n9819) );
  BUF_X1 U341 ( .A(n9232), .Z(n9818) );
  BUF_X1 U342 ( .A(n9232), .Z(n9817) );
  BUF_X1 U343 ( .A(n9232), .Z(n9816) );
  BUF_X1 U344 ( .A(n9232), .Z(n9815) );
  BUF_X1 U345 ( .A(n9232), .Z(n9814) );
  BUF_X1 U346 ( .A(n9227), .Z(n9693) );
  BUF_X1 U347 ( .A(n9227), .Z(n9694) );
  BUF_X1 U348 ( .A(n9227), .Z(n9695) );
  BUF_X1 U349 ( .A(n9227), .Z(n9696) );
  BUF_X1 U350 ( .A(n9227), .Z(n9697) );
  BUF_X1 U351 ( .A(n9227), .Z(n9698) );
  BUF_X1 U352 ( .A(n9696), .Z(n9699) );
  BUF_X1 U353 ( .A(n9697), .Z(n9700) );
  BUF_X1 U354 ( .A(n9805), .Z(n9810) );
  BUF_X1 U355 ( .A(n9804), .Z(n9809) );
  BUF_X1 U356 ( .A(n9236), .Z(n9808) );
  BUF_X1 U357 ( .A(n9236), .Z(n9807) );
  BUF_X1 U358 ( .A(n9236), .Z(n9806) );
  BUF_X1 U359 ( .A(n9236), .Z(n9805) );
  BUF_X1 U360 ( .A(n9236), .Z(n9804) );
  BUF_X1 U361 ( .A(n9236), .Z(n9803) );
  BUF_X1 U362 ( .A(n9673), .Z(n9678) );
  BUF_X1 U363 ( .A(n9672), .Z(n9677) );
  BUF_X1 U364 ( .A(n9230), .Z(n9676) );
  BUF_X1 U365 ( .A(n9230), .Z(n9675) );
  BUF_X1 U366 ( .A(n9230), .Z(n9674) );
  BUF_X1 U367 ( .A(n9230), .Z(n9673) );
  BUF_X1 U368 ( .A(n9230), .Z(n9672) );
  BUF_X1 U369 ( .A(n9230), .Z(n9671) );
  BUF_X1 U370 ( .A(n9794), .Z(n9799) );
  BUF_X1 U371 ( .A(n9793), .Z(n9798) );
  BUF_X1 U372 ( .A(n9237), .Z(n9797) );
  BUF_X1 U373 ( .A(n9237), .Z(n9796) );
  BUF_X1 U374 ( .A(n9237), .Z(n9795) );
  BUF_X1 U375 ( .A(n9237), .Z(n9794) );
  BUF_X1 U376 ( .A(n9237), .Z(n9793) );
  BUF_X1 U377 ( .A(n9237), .Z(n9792) );
  BUF_X1 U378 ( .A(n9884), .Z(n9880) );
  BUF_X1 U379 ( .A(n9884), .Z(n9882) );
  BUF_X1 U380 ( .A(n9884), .Z(n9881) );
  BUF_X1 U381 ( .A(n1516), .Z(n9364) );
  BUF_X1 U382 ( .A(n1526), .Z(n9340) );
  BUF_X1 U383 ( .A(n1516), .Z(n9365) );
  BUF_X1 U384 ( .A(n1526), .Z(n9341) );
  BUF_X1 U385 ( .A(n872), .Z(n9508) );
  BUF_X1 U386 ( .A(n872), .Z(n9509) );
  BUF_X1 U387 ( .A(n877), .Z(n9496) );
  BUF_X1 U388 ( .A(n901), .Z(n9448) );
  BUF_X1 U389 ( .A(n906), .Z(n9436) );
  BUF_X1 U390 ( .A(n882), .Z(n9484) );
  BUF_X1 U391 ( .A(n906), .Z(n9437) );
  BUF_X1 U392 ( .A(n877), .Z(n9497) );
  BUF_X1 U393 ( .A(n867), .Z(n9521) );
  BUF_X1 U394 ( .A(n901), .Z(n9449) );
  BUF_X1 U395 ( .A(n882), .Z(n9485) );
  BUF_X1 U396 ( .A(n1487), .Z(n9424) );
  BUF_X1 U397 ( .A(n1492), .Z(n9412) );
  BUF_X1 U398 ( .A(n1497), .Z(n9400) );
  BUF_X1 U399 ( .A(n1502), .Z(n9388) );
  BUF_X1 U400 ( .A(n1511), .Z(n9376) );
  BUF_X1 U401 ( .A(n1521), .Z(n9352) );
  BUF_X1 U402 ( .A(n1487), .Z(n9425) );
  BUF_X1 U403 ( .A(n1492), .Z(n9413) );
  BUF_X1 U404 ( .A(n1497), .Z(n9401) );
  BUF_X1 U405 ( .A(n1502), .Z(n9389) );
  BUF_X1 U406 ( .A(n1511), .Z(n9377) );
  BUF_X1 U407 ( .A(n1521), .Z(n9353) );
  BUF_X1 U408 ( .A(n893), .Z(n9469) );
  BUF_X1 U409 ( .A(n874), .Z(n9505) );
  BUF_X1 U410 ( .A(n898), .Z(n9457) );
  BUF_X1 U411 ( .A(n884), .Z(n9481) );
  BUF_X1 U412 ( .A(n903), .Z(n9445) );
  BUF_X1 U413 ( .A(n908), .Z(n9433) );
  BUF_X1 U414 ( .A(n879), .Z(n9493) );
  BUF_X1 U415 ( .A(n874), .Z(n9506) );
  BUF_X1 U416 ( .A(n893), .Z(n9470) );
  BUF_X1 U417 ( .A(n898), .Z(n9458) );
  BUF_X1 U418 ( .A(n903), .Z(n9446) );
  BUF_X1 U419 ( .A(n869), .Z(n9518) );
  BUF_X1 U420 ( .A(n884), .Z(n9482) );
  BUF_X1 U421 ( .A(n879), .Z(n9494) );
  BUF_X1 U422 ( .A(n908), .Z(n9434) );
  BUF_X1 U423 ( .A(n1489), .Z(n9421) );
  BUF_X1 U424 ( .A(n1494), .Z(n9409) );
  BUF_X1 U425 ( .A(n1499), .Z(n9397) );
  BUF_X1 U426 ( .A(n1504), .Z(n9385) );
  BUF_X1 U427 ( .A(n1513), .Z(n9373) );
  BUF_X1 U428 ( .A(n1523), .Z(n9349) );
  BUF_X1 U429 ( .A(n1518), .Z(n9361) );
  BUF_X1 U430 ( .A(n1528), .Z(n9337) );
  BUF_X1 U431 ( .A(n1489), .Z(n9422) );
  BUF_X1 U432 ( .A(n1494), .Z(n9410) );
  BUF_X1 U433 ( .A(n1499), .Z(n9398) );
  BUF_X1 U434 ( .A(n1504), .Z(n9386) );
  BUF_X1 U435 ( .A(n1513), .Z(n9374) );
  BUF_X1 U436 ( .A(n1523), .Z(n9350) );
  BUF_X1 U437 ( .A(n1518), .Z(n9362) );
  BUF_X1 U438 ( .A(n1528), .Z(n9338) );
  BUF_X1 U439 ( .A(n905), .Z(n9439) );
  BUF_X1 U440 ( .A(n905), .Z(n9440) );
  BUF_X1 U441 ( .A(n1515), .Z(n9367) );
  BUF_X1 U442 ( .A(n1525), .Z(n9343) );
  BUF_X1 U443 ( .A(n1515), .Z(n9368) );
  BUF_X1 U444 ( .A(n1525), .Z(n9344) );
  BUF_X1 U445 ( .A(n871), .Z(n9511) );
  BUF_X1 U446 ( .A(n871), .Z(n9512) );
  BUF_X1 U447 ( .A(n1491), .Z(n9415) );
  BUF_X1 U448 ( .A(n1491), .Z(n9416) );
  BUF_X1 U449 ( .A(n900), .Z(n9451) );
  BUF_X1 U450 ( .A(n876), .Z(n9499) );
  BUF_X1 U451 ( .A(n881), .Z(n9487) );
  BUF_X1 U452 ( .A(n866), .Z(n9524) );
  BUF_X1 U453 ( .A(n900), .Z(n9452) );
  BUF_X1 U454 ( .A(n876), .Z(n9500) );
  BUF_X1 U455 ( .A(n881), .Z(n9488) );
  BUF_X1 U456 ( .A(n1486), .Z(n9427) );
  BUF_X1 U457 ( .A(n1496), .Z(n9403) );
  BUF_X1 U458 ( .A(n1501), .Z(n9391) );
  BUF_X1 U459 ( .A(n1510), .Z(n9379) );
  BUF_X1 U460 ( .A(n1520), .Z(n9355) );
  BUF_X1 U461 ( .A(n1486), .Z(n9428) );
  BUF_X1 U462 ( .A(n1496), .Z(n9404) );
  BUF_X1 U463 ( .A(n1501), .Z(n9392) );
  BUF_X1 U464 ( .A(n1510), .Z(n9380) );
  BUF_X1 U465 ( .A(n1520), .Z(n9356) );
  BUF_X1 U466 ( .A(n867), .Z(n9520) );
  BUF_X1 U467 ( .A(n869), .Z(n9517) );
  BUF_X1 U468 ( .A(n866), .Z(n9523) );
  BUF_X1 U469 ( .A(n885), .Z(n9478) );
  BUF_X1 U470 ( .A(n894), .Z(n9466) );
  BUF_X1 U471 ( .A(n870), .Z(n9514) );
  BUF_X1 U472 ( .A(n899), .Z(n9454) );
  BUF_X1 U473 ( .A(n880), .Z(n9490) );
  BUF_X1 U474 ( .A(n875), .Z(n9502) );
  BUF_X1 U475 ( .A(n904), .Z(n9442) );
  BUF_X1 U476 ( .A(n875), .Z(n9503) );
  BUF_X1 U477 ( .A(n870), .Z(n9515) );
  BUF_X1 U478 ( .A(n894), .Z(n9467) );
  BUF_X1 U479 ( .A(n899), .Z(n9455) );
  BUF_X1 U480 ( .A(n885), .Z(n9479) );
  BUF_X1 U481 ( .A(n880), .Z(n9491) );
  BUF_X1 U482 ( .A(n904), .Z(n9443) );
  BUF_X1 U483 ( .A(n909), .Z(n9430) );
  BUF_X1 U484 ( .A(n909), .Z(n9431) );
  BUF_X1 U485 ( .A(n1490), .Z(n9419) );
  BUF_X1 U486 ( .A(n1495), .Z(n9407) );
  BUF_X1 U487 ( .A(n1500), .Z(n9395) );
  BUF_X1 U488 ( .A(n1505), .Z(n9383) );
  BUF_X1 U489 ( .A(n1514), .Z(n9371) );
  BUF_X1 U490 ( .A(n1524), .Z(n9347) );
  BUF_X1 U491 ( .A(n1519), .Z(n9359) );
  BUF_X1 U492 ( .A(n1529), .Z(n9335) );
  BUF_X1 U493 ( .A(n1490), .Z(n9418) );
  BUF_X1 U494 ( .A(n1495), .Z(n9406) );
  BUF_X1 U495 ( .A(n1500), .Z(n9394) );
  BUF_X1 U496 ( .A(n1505), .Z(n9382) );
  BUF_X1 U497 ( .A(n1514), .Z(n9370) );
  BUF_X1 U498 ( .A(n1524), .Z(n9346) );
  BUF_X1 U499 ( .A(n1519), .Z(n9358) );
  BUF_X1 U500 ( .A(n1529), .Z(n9334) );
  BUF_X1 U501 ( .A(n891), .Z(n9472) );
  BUF_X1 U502 ( .A(n896), .Z(n9460) );
  BUF_X1 U503 ( .A(n896), .Z(n9461) );
  BUF_X1 U504 ( .A(n891), .Z(n9473) );
  BUF_X1 U505 ( .A(n1516), .Z(n9366) );
  BUF_X1 U506 ( .A(n1526), .Z(n9342) );
  BUF_X1 U507 ( .A(n1492), .Z(n9414) );
  BUF_X1 U508 ( .A(n882), .Z(n9486) );
  BUF_X1 U509 ( .A(n867), .Z(n9522) );
  BUF_X1 U510 ( .A(n877), .Z(n9498) );
  BUF_X1 U511 ( .A(n896), .Z(n9462) );
  BUF_X1 U512 ( .A(n891), .Z(n9474) );
  BUF_X1 U513 ( .A(n901), .Z(n9450) );
  BUF_X1 U514 ( .A(n872), .Z(n9510) );
  BUF_X1 U515 ( .A(n906), .Z(n9438) );
  BUF_X1 U516 ( .A(n1487), .Z(n9426) );
  BUF_X1 U517 ( .A(n1497), .Z(n9402) );
  BUF_X1 U518 ( .A(n1502), .Z(n9390) );
  BUF_X1 U519 ( .A(n1511), .Z(n9378) );
  BUF_X1 U520 ( .A(n1521), .Z(n9354) );
  BUF_X1 U521 ( .A(n890), .Z(n9475) );
  BUF_X1 U522 ( .A(n895), .Z(n9463) );
  BUF_X1 U523 ( .A(n890), .Z(n9476) );
  BUF_X1 U524 ( .A(n895), .Z(n9464) );
  BUF_X1 U525 ( .A(n898), .Z(n9459) );
  BUF_X1 U526 ( .A(n869), .Z(n9519) );
  BUF_X1 U527 ( .A(n893), .Z(n9471) );
  BUF_X1 U528 ( .A(n884), .Z(n9483) );
  BUF_X1 U529 ( .A(n903), .Z(n9447) );
  BUF_X1 U530 ( .A(n874), .Z(n9507) );
  BUF_X1 U531 ( .A(n879), .Z(n9495) );
  BUF_X1 U532 ( .A(n908), .Z(n9435) );
  BUF_X1 U533 ( .A(n1489), .Z(n9423) );
  BUF_X1 U534 ( .A(n1494), .Z(n9411) );
  BUF_X1 U535 ( .A(n1499), .Z(n9399) );
  BUF_X1 U536 ( .A(n1504), .Z(n9387) );
  BUF_X1 U537 ( .A(n1513), .Z(n9375) );
  BUF_X1 U538 ( .A(n1523), .Z(n9351) );
  BUF_X1 U539 ( .A(n1518), .Z(n9363) );
  BUF_X1 U540 ( .A(n1528), .Z(n9339) );
  BUF_X1 U541 ( .A(n905), .Z(n9441) );
  BUF_X1 U542 ( .A(n1515), .Z(n9369) );
  BUF_X1 U543 ( .A(n1525), .Z(n9345) );
  BUF_X1 U544 ( .A(n1491), .Z(n9417) );
  BUF_X1 U545 ( .A(n881), .Z(n9489) );
  BUF_X1 U546 ( .A(n890), .Z(n9477) );
  BUF_X1 U547 ( .A(n866), .Z(n9525) );
  BUF_X1 U548 ( .A(n895), .Z(n9465) );
  BUF_X1 U549 ( .A(n871), .Z(n9513) );
  BUF_X1 U550 ( .A(n900), .Z(n9453) );
  BUF_X1 U551 ( .A(n876), .Z(n9501) );
  BUF_X1 U552 ( .A(n1486), .Z(n9429) );
  BUF_X1 U553 ( .A(n1496), .Z(n9405) );
  BUF_X1 U554 ( .A(n1501), .Z(n9393) );
  BUF_X1 U555 ( .A(n1510), .Z(n9381) );
  BUF_X1 U556 ( .A(n1520), .Z(n9357) );
  BUF_X1 U557 ( .A(n875), .Z(n9504) );
  BUF_X1 U558 ( .A(n885), .Z(n9480) );
  BUF_X1 U559 ( .A(n899), .Z(n9456) );
  BUF_X1 U560 ( .A(n909), .Z(n9432) );
  BUF_X1 U561 ( .A(n894), .Z(n9468) );
  BUF_X1 U562 ( .A(n880), .Z(n9492) );
  BUF_X1 U563 ( .A(n904), .Z(n9444) );
  BUF_X1 U564 ( .A(n1514), .Z(n9372) );
  BUF_X1 U565 ( .A(n1524), .Z(n9348) );
  BUF_X1 U566 ( .A(n1519), .Z(n9360) );
  BUF_X1 U567 ( .A(n1529), .Z(n9336) );
  BUF_X1 U568 ( .A(n1490), .Z(n9420) );
  BUF_X1 U569 ( .A(n1495), .Z(n9408) );
  BUF_X1 U570 ( .A(n1500), .Z(n9396) );
  BUF_X1 U571 ( .A(n1505), .Z(n9384) );
  BUF_X1 U572 ( .A(n870), .Z(n9516) );
  BUF_X1 U573 ( .A(n815), .Z(n9874) );
  BUF_X1 U574 ( .A(n815), .Z(n9873) );
  BUF_X1 U575 ( .A(n815), .Z(n9872) );
  BUF_X1 U576 ( .A(n815), .Z(n9871) );
  BUF_X1 U577 ( .A(n815), .Z(n9870) );
  BUF_X1 U578 ( .A(n815), .Z(n9869) );
  BUF_X1 U579 ( .A(n815), .Z(n9875) );
  INV_X1 U580 ( .A(n9876), .ZN(n9884) );
  NOR3_X1 U581 ( .A1(n9920), .A2(n9919), .A3(n9921), .ZN(n824) );
  AND3_X1 U582 ( .A1(n9918), .A2(n9917), .A3(n849), .ZN(n830) );
  BUF_X1 U583 ( .A(n9916), .Z(n9331) );
  BUF_X1 U584 ( .A(n9915), .Z(n9328) );
  BUF_X1 U585 ( .A(n9914), .Z(n9325) );
  BUF_X1 U586 ( .A(n9913), .Z(n9322) );
  BUF_X1 U587 ( .A(n9912), .Z(n9319) );
  BUF_X1 U588 ( .A(n9911), .Z(n9316) );
  BUF_X1 U589 ( .A(n9910), .Z(n9313) );
  BUF_X1 U590 ( .A(n9909), .Z(n9310) );
  BUF_X1 U591 ( .A(n9908), .Z(n9307) );
  BUF_X1 U592 ( .A(n9907), .Z(n9304) );
  BUF_X1 U593 ( .A(n9906), .Z(n9301) );
  BUF_X1 U594 ( .A(n9905), .Z(n9298) );
  BUF_X1 U595 ( .A(n9904), .Z(n9295) );
  BUF_X1 U596 ( .A(n9903), .Z(n9292) );
  BUF_X1 U597 ( .A(n9902), .Z(n9289) );
  BUF_X1 U598 ( .A(n9901), .Z(n9286) );
  BUF_X1 U599 ( .A(n9900), .Z(n9283) );
  BUF_X1 U600 ( .A(n9899), .Z(n9280) );
  BUF_X1 U601 ( .A(n9898), .Z(n9277) );
  BUF_X1 U602 ( .A(n9897), .Z(n9274) );
  BUF_X1 U603 ( .A(n9896), .Z(n9271) );
  BUF_X1 U604 ( .A(n9895), .Z(n9268) );
  BUF_X1 U605 ( .A(n9894), .Z(n9265) );
  BUF_X1 U606 ( .A(n9893), .Z(n9262) );
  BUF_X1 U607 ( .A(n9892), .Z(n9259) );
  BUF_X1 U608 ( .A(n9891), .Z(n9256) );
  BUF_X1 U609 ( .A(n9890), .Z(n9253) );
  BUF_X1 U610 ( .A(n9889), .Z(n9250) );
  BUF_X1 U611 ( .A(n9888), .Z(n9247) );
  BUF_X1 U612 ( .A(n9887), .Z(n9244) );
  BUF_X1 U613 ( .A(n9886), .Z(n9241) );
  BUF_X1 U614 ( .A(n9885), .Z(n9238) );
  BUF_X1 U615 ( .A(n9916), .Z(n9332) );
  BUF_X1 U616 ( .A(n9915), .Z(n9329) );
  BUF_X1 U617 ( .A(n9914), .Z(n9326) );
  BUF_X1 U618 ( .A(n9913), .Z(n9323) );
  BUF_X1 U619 ( .A(n9912), .Z(n9320) );
  BUF_X1 U620 ( .A(n9911), .Z(n9317) );
  BUF_X1 U621 ( .A(n9910), .Z(n9314) );
  BUF_X1 U622 ( .A(n9909), .Z(n9311) );
  BUF_X1 U623 ( .A(n9908), .Z(n9308) );
  BUF_X1 U624 ( .A(n9907), .Z(n9305) );
  BUF_X1 U625 ( .A(n9906), .Z(n9302) );
  BUF_X1 U626 ( .A(n9905), .Z(n9299) );
  BUF_X1 U627 ( .A(n9904), .Z(n9296) );
  BUF_X1 U628 ( .A(n9903), .Z(n9293) );
  BUF_X1 U629 ( .A(n9902), .Z(n9290) );
  BUF_X1 U630 ( .A(n9901), .Z(n9287) );
  BUF_X1 U631 ( .A(n9900), .Z(n9284) );
  BUF_X1 U632 ( .A(n9899), .Z(n9281) );
  BUF_X1 U633 ( .A(n9898), .Z(n9278) );
  BUF_X1 U634 ( .A(n9897), .Z(n9275) );
  BUF_X1 U635 ( .A(n9896), .Z(n9272) );
  BUF_X1 U636 ( .A(n9895), .Z(n9269) );
  BUF_X1 U637 ( .A(n9894), .Z(n9266) );
  BUF_X1 U638 ( .A(n9893), .Z(n9263) );
  BUF_X1 U639 ( .A(n9892), .Z(n9260) );
  BUF_X1 U640 ( .A(n9891), .Z(n9257) );
  BUF_X1 U641 ( .A(n9890), .Z(n9254) );
  BUF_X1 U642 ( .A(n9889), .Z(n9251) );
  BUF_X1 U643 ( .A(n9888), .Z(n9248) );
  BUF_X1 U644 ( .A(n9887), .Z(n9245) );
  BUF_X1 U645 ( .A(n9886), .Z(n9242) );
  BUF_X1 U646 ( .A(n9885), .Z(n9239) );
  NAND2_X1 U647 ( .A1(n1459), .A2(n1458), .ZN(n866) );
  NAND2_X1 U648 ( .A1(n1457), .A2(n1470), .ZN(n896) );
  AOI22_X1 U649 ( .A1(n9483), .A2(n10194), .B1(n9478), .B2(n10554), .ZN(n883)
         );
  AOI22_X1 U650 ( .A1(n9483), .A2(n10200), .B1(n9478), .B2(n10560), .ZN(n1009)
         );
  AOI22_X1 U651 ( .A1(n9483), .A2(n10197), .B1(n9478), .B2(n10557), .ZN(n955)
         );
  AOI22_X1 U652 ( .A1(n9483), .A2(n10201), .B1(n9478), .B2(n10561), .ZN(n1027)
         );
  AOI22_X1 U653 ( .A1(n9483), .A2(n10196), .B1(n9478), .B2(n10556), .ZN(n937)
         );
  AOI22_X1 U654 ( .A1(n9483), .A2(n10199), .B1(n9478), .B2(n10559), .ZN(n991)
         );
  AOI22_X1 U655 ( .A1(n9483), .A2(n10195), .B1(n9478), .B2(n10555), .ZN(n919)
         );
  AOI22_X1 U656 ( .A1(n9483), .A2(n10198), .B1(n9478), .B2(n10558), .ZN(n973)
         );
  NAND2_X1 U657 ( .A1(n2084), .A2(n2088), .ZN(n1501) );
  NAND2_X1 U658 ( .A1(n2083), .A2(n2088), .ZN(n1502) );
  NAND2_X1 U659 ( .A1(n1477), .A2(n1459), .ZN(n905) );
  NAND2_X1 U660 ( .A1(n1461), .A2(n1460), .ZN(n872) );
  NAND2_X1 U661 ( .A1(n1461), .A2(n1458), .ZN(n867) );
  NAND2_X1 U662 ( .A1(n816), .A2(n817), .ZN(n815) );
  BUF_X1 U663 ( .A(n9916), .Z(n9333) );
  BUF_X1 U664 ( .A(n9915), .Z(n9330) );
  BUF_X1 U665 ( .A(n9914), .Z(n9327) );
  BUF_X1 U666 ( .A(n9913), .Z(n9324) );
  BUF_X1 U667 ( .A(n9912), .Z(n9321) );
  BUF_X1 U668 ( .A(n9911), .Z(n9318) );
  BUF_X1 U669 ( .A(n9910), .Z(n9315) );
  BUF_X1 U670 ( .A(n9909), .Z(n9312) );
  BUF_X1 U671 ( .A(n9908), .Z(n9309) );
  BUF_X1 U672 ( .A(n9907), .Z(n9306) );
  BUF_X1 U673 ( .A(n9906), .Z(n9303) );
  BUF_X1 U674 ( .A(n9905), .Z(n9300) );
  BUF_X1 U675 ( .A(n9904), .Z(n9297) );
  BUF_X1 U676 ( .A(n9903), .Z(n9294) );
  BUF_X1 U677 ( .A(n9902), .Z(n9291) );
  BUF_X1 U678 ( .A(n9901), .Z(n9288) );
  BUF_X1 U679 ( .A(n9900), .Z(n9285) );
  BUF_X1 U680 ( .A(n9899), .Z(n9282) );
  BUF_X1 U681 ( .A(n9898), .Z(n9279) );
  BUF_X1 U682 ( .A(n9897), .Z(n9276) );
  BUF_X1 U683 ( .A(n9896), .Z(n9273) );
  BUF_X1 U684 ( .A(n9895), .Z(n9270) );
  BUF_X1 U685 ( .A(n9894), .Z(n9267) );
  BUF_X1 U686 ( .A(n9893), .Z(n9264) );
  BUF_X1 U687 ( .A(n9892), .Z(n9261) );
  BUF_X1 U688 ( .A(n9891), .Z(n9258) );
  BUF_X1 U689 ( .A(n9890), .Z(n9255) );
  BUF_X1 U690 ( .A(n9889), .Z(n9252) );
  BUF_X1 U691 ( .A(n9888), .Z(n9249) );
  BUF_X1 U692 ( .A(n9887), .Z(n9246) );
  BUF_X1 U693 ( .A(n9886), .Z(n9243) );
  BUF_X1 U694 ( .A(n9885), .Z(n9240) );
  NAND2_X1 U695 ( .A1(n2095), .A2(n2084), .ZN(n1515) );
  NAND2_X1 U696 ( .A1(n2095), .A2(n2083), .ZN(n1516) );
  NAND2_X1 U697 ( .A1(n2098), .A2(n2084), .ZN(n1525) );
  NAND2_X1 U698 ( .A1(n2098), .A2(n2083), .ZN(n1526) );
  NAND2_X1 U699 ( .A1(n1477), .A2(n1461), .ZN(n906) );
  NAND2_X1 U700 ( .A1(n1464), .A2(n1460), .ZN(n881) );
  NAND2_X1 U701 ( .A1(n2077), .A2(n2085), .ZN(n1492) );
  NAND2_X1 U702 ( .A1(n2077), .A2(n2086), .ZN(n1491) );
  NAND2_X1 U703 ( .A1(n1458), .A2(n1464), .ZN(n871) );
  NAND2_X1 U704 ( .A1(n1470), .A2(n1464), .ZN(n891) );
  NAND2_X1 U705 ( .A1(n1477), .A2(n1464), .ZN(n895) );
  NAND2_X1 U706 ( .A1(n1468), .A2(n1470), .ZN(n890) );
  AND2_X1 U707 ( .A1(n1459), .A2(n1470), .ZN(n898) );
  AND2_X1 U708 ( .A1(n1459), .A2(n1460), .ZN(n869) );
  NAND2_X1 U709 ( .A1(n1458), .A2(n1468), .ZN(n877) );
  NAND2_X1 U710 ( .A1(n1477), .A2(n1468), .ZN(n901) );
  NAND2_X1 U711 ( .A1(n1458), .A2(n1467), .ZN(n876) );
  NAND2_X1 U712 ( .A1(n2079), .A2(n2088), .ZN(n1496) );
  NAND2_X1 U713 ( .A1(n2078), .A2(n2088), .ZN(n1497) );
  AND2_X1 U714 ( .A1(n1457), .A2(n1460), .ZN(n875) );
  AND2_X1 U715 ( .A1(n1457), .A2(n1458), .ZN(n870) );
  NAND2_X1 U716 ( .A1(n1466), .A2(n1460), .ZN(n882) );
  NAND2_X1 U717 ( .A1(n2095), .A2(n2079), .ZN(n1510) );
  NAND2_X1 U718 ( .A1(n2095), .A2(n2078), .ZN(n1511) );
  NAND2_X1 U719 ( .A1(n2098), .A2(n2079), .ZN(n1520) );
  NAND2_X1 U720 ( .A1(n2098), .A2(n2078), .ZN(n1521) );
  NAND2_X1 U721 ( .A1(n1477), .A2(n1467), .ZN(n900) );
  NAND2_X1 U722 ( .A1(n2077), .A2(n2081), .ZN(n1486) );
  NAND2_X1 U723 ( .A1(n2077), .A2(n2080), .ZN(n1487) );
  AND2_X1 U724 ( .A1(n1477), .A2(n1457), .ZN(n909) );
  AND2_X1 U725 ( .A1(n1461), .A2(n1470), .ZN(n899) );
  AND2_X1 U726 ( .A1(n2085), .A2(n2088), .ZN(n1505) );
  AND2_X1 U727 ( .A1(n2086), .A2(n2088), .ZN(n1504) );
  AND2_X1 U728 ( .A1(n2077), .A2(n2083), .ZN(n1495) );
  AND2_X1 U729 ( .A1(n2077), .A2(n2084), .ZN(n1494) );
  AND2_X1 U730 ( .A1(n1463), .A2(n1470), .ZN(n893) );
  AND2_X1 U731 ( .A1(n1463), .A2(n1460), .ZN(n874) );
  AND2_X1 U732 ( .A1(n1463), .A2(n1458), .ZN(n908) );
  AND2_X1 U733 ( .A1(n2095), .A2(n2085), .ZN(n1519) );
  AND2_X1 U734 ( .A1(n2095), .A2(n2086), .ZN(n1518) );
  AND2_X1 U735 ( .A1(n2098), .A2(n2085), .ZN(n1529) );
  AND2_X1 U736 ( .A1(n2098), .A2(n2086), .ZN(n1528) );
  AND2_X1 U737 ( .A1(n1477), .A2(n1463), .ZN(n903) );
  AND2_X1 U738 ( .A1(n1468), .A2(n1460), .ZN(n885) );
  AND2_X1 U739 ( .A1(n1458), .A2(n1466), .ZN(n880) );
  AND2_X1 U740 ( .A1(n1477), .A2(n1466), .ZN(n904) );
  AND2_X1 U741 ( .A1(n2077), .A2(n2079), .ZN(n1489) );
  AND2_X1 U742 ( .A1(n2077), .A2(n2078), .ZN(n1490) );
  AND2_X1 U743 ( .A1(n2095), .A2(n2081), .ZN(n1513) );
  AND2_X1 U744 ( .A1(n2095), .A2(n2080), .ZN(n1514) );
  AND2_X1 U745 ( .A1(n2098), .A2(n2081), .ZN(n1523) );
  AND2_X1 U746 ( .A1(n2098), .A2(n2080), .ZN(n1524) );
  AND2_X1 U747 ( .A1(n1470), .A2(n1466), .ZN(n884) );
  AND2_X1 U748 ( .A1(n2081), .A2(n2088), .ZN(n1499) );
  AND2_X1 U749 ( .A1(n2080), .A2(n2088), .ZN(n1500) );
  AND2_X1 U750 ( .A1(n1467), .A2(n1460), .ZN(n879) );
  AND2_X1 U751 ( .A1(n1467), .A2(n1470), .ZN(n894) );
  NOR3_X1 U752 ( .A1(ADD_WR[0]), .A2(ADD_WR[1]), .A3(n9919), .ZN(n817) );
  NOR3_X1 U753 ( .A1(ADD_WR[0]), .A2(ADD_WR[2]), .A3(n9920), .ZN(n822) );
  NOR3_X1 U754 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n819) );
  NOR3_X1 U755 ( .A1(n9919), .A2(ADD_WR[1]), .A3(n9921), .ZN(n827) );
  NOR3_X1 U756 ( .A1(n9919), .A2(ADD_WR[0]), .A3(n9920), .ZN(n847) );
  NOR3_X1 U757 ( .A1(n9920), .A2(ADD_WR[2]), .A3(n9921), .ZN(n845) );
  NOR3_X1 U758 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(n9921), .ZN(n842) );
  NOR3_X1 U759 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[2]), .A3(n10663), .ZN(n2084) );
  NOR3_X1 U760 ( .A1(n10664), .A2(ADD_RD2[2]), .A3(n10663), .ZN(n2083) );
  NOR3_X1 U761 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[2]), .A3(n10659), .ZN(n1461) );
  NOR3_X1 U762 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n10664), .ZN(n2085) );
  NOR3_X1 U763 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(ADD_RD2[0]), .ZN(n2086)
         );
  NOR3_X1 U764 ( .A1(n10660), .A2(ADD_RD1[2]), .A3(n10659), .ZN(n1463) );
  NOR4_X1 U765 ( .A1(n1928), .A2(n1929), .A3(n1930), .A4(n1931), .ZN(n1927) );
  OAI221_X1 U766 ( .B1(n8574), .B2(n9391), .C1(n8550), .C2(n9388), .A(n1935), 
        .ZN(n1928) );
  OAI221_X1 U767 ( .B1(n8486), .B2(n9403), .C1(n8247), .C2(n9400), .A(n1934), 
        .ZN(n1929) );
  OAI221_X1 U768 ( .B1(n8447), .B2(n9415), .C1(n8415), .C2(n9412), .A(n1933), 
        .ZN(n1930) );
  NOR4_X1 U769 ( .A1(n1910), .A2(n1911), .A3(n1912), .A4(n1913), .ZN(n1909) );
  OAI221_X1 U770 ( .B1(n8575), .B2(n9391), .C1(n8551), .C2(n9388), .A(n1917), 
        .ZN(n1910) );
  OAI221_X1 U771 ( .B1(n8487), .B2(n9403), .C1(n8248), .C2(n9400), .A(n1916), 
        .ZN(n1911) );
  OAI221_X1 U772 ( .B1(n8448), .B2(n9415), .C1(n8416), .C2(n9412), .A(n1915), 
        .ZN(n1912) );
  NOR4_X1 U773 ( .A1(n1892), .A2(n1893), .A3(n1894), .A4(n1895), .ZN(n1891) );
  OAI221_X1 U774 ( .B1(n8576), .B2(n9391), .C1(n8552), .C2(n9388), .A(n1899), 
        .ZN(n1892) );
  OAI221_X1 U775 ( .B1(n8488), .B2(n9403), .C1(n8249), .C2(n9400), .A(n1898), 
        .ZN(n1893) );
  OAI221_X1 U776 ( .B1(n8449), .B2(n9415), .C1(n8417), .C2(n9412), .A(n1897), 
        .ZN(n1894) );
  NOR4_X1 U777 ( .A1(n1874), .A2(n1875), .A3(n1876), .A4(n1877), .ZN(n1873) );
  OAI221_X1 U778 ( .B1(n8577), .B2(n9391), .C1(n8553), .C2(n9388), .A(n1881), 
        .ZN(n1874) );
  OAI221_X1 U779 ( .B1(n8489), .B2(n9403), .C1(n8250), .C2(n9400), .A(n1880), 
        .ZN(n1875) );
  OAI221_X1 U780 ( .B1(n8450), .B2(n9415), .C1(n8418), .C2(n9412), .A(n1879), 
        .ZN(n1876) );
  NOR4_X1 U781 ( .A1(n1856), .A2(n1857), .A3(n1858), .A4(n1859), .ZN(n1855) );
  OAI221_X1 U782 ( .B1(n8578), .B2(n9392), .C1(n8554), .C2(n9389), .A(n1863), 
        .ZN(n1856) );
  OAI221_X1 U783 ( .B1(n8490), .B2(n9404), .C1(n8251), .C2(n9401), .A(n1862), 
        .ZN(n1857) );
  OAI221_X1 U784 ( .B1(n8451), .B2(n9416), .C1(n8419), .C2(n9413), .A(n1861), 
        .ZN(n1858) );
  NOR4_X1 U785 ( .A1(n1838), .A2(n1839), .A3(n1840), .A4(n1841), .ZN(n1837) );
  OAI221_X1 U786 ( .B1(n8579), .B2(n9392), .C1(n8555), .C2(n9389), .A(n1845), 
        .ZN(n1838) );
  OAI221_X1 U787 ( .B1(n8491), .B2(n9404), .C1(n8252), .C2(n9401), .A(n1844), 
        .ZN(n1839) );
  OAI221_X1 U788 ( .B1(n8452), .B2(n9416), .C1(n8420), .C2(n9413), .A(n1843), 
        .ZN(n1840) );
  NOR4_X1 U789 ( .A1(n1820), .A2(n1821), .A3(n1822), .A4(n1823), .ZN(n1819) );
  OAI221_X1 U790 ( .B1(n8580), .B2(n9392), .C1(n8556), .C2(n9389), .A(n1827), 
        .ZN(n1820) );
  OAI221_X1 U791 ( .B1(n8492), .B2(n9404), .C1(n8253), .C2(n9401), .A(n1826), 
        .ZN(n1821) );
  OAI221_X1 U792 ( .B1(n8453), .B2(n9416), .C1(n8421), .C2(n9413), .A(n1825), 
        .ZN(n1822) );
  NOR4_X1 U793 ( .A1(n1802), .A2(n1803), .A3(n1804), .A4(n1805), .ZN(n1801) );
  OAI221_X1 U794 ( .B1(n8581), .B2(n9392), .C1(n8557), .C2(n9389), .A(n1809), 
        .ZN(n1802) );
  OAI221_X1 U795 ( .B1(n8493), .B2(n9404), .C1(n8254), .C2(n9401), .A(n1808), 
        .ZN(n1803) );
  OAI221_X1 U796 ( .B1(n8454), .B2(n9416), .C1(n8422), .C2(n9413), .A(n1807), 
        .ZN(n1804) );
  NOR4_X1 U797 ( .A1(n1784), .A2(n1785), .A3(n1786), .A4(n1787), .ZN(n1783) );
  OAI221_X1 U798 ( .B1(n8582), .B2(n9392), .C1(n8558), .C2(n9389), .A(n1791), 
        .ZN(n1784) );
  OAI221_X1 U799 ( .B1(n8494), .B2(n9404), .C1(n8255), .C2(n9401), .A(n1790), 
        .ZN(n1785) );
  OAI221_X1 U800 ( .B1(n8455), .B2(n9416), .C1(n8423), .C2(n9413), .A(n1789), 
        .ZN(n1786) );
  NOR4_X1 U801 ( .A1(n1766), .A2(n1767), .A3(n1768), .A4(n1769), .ZN(n1765) );
  OAI221_X1 U802 ( .B1(n8583), .B2(n9392), .C1(n8559), .C2(n9389), .A(n1773), 
        .ZN(n1766) );
  OAI221_X1 U803 ( .B1(n8495), .B2(n9404), .C1(n8256), .C2(n9401), .A(n1772), 
        .ZN(n1767) );
  OAI221_X1 U804 ( .B1(n8456), .B2(n9416), .C1(n8424), .C2(n9413), .A(n1771), 
        .ZN(n1768) );
  NOR4_X1 U805 ( .A1(n1748), .A2(n1749), .A3(n1750), .A4(n1751), .ZN(n1747) );
  OAI221_X1 U806 ( .B1(n8584), .B2(n9392), .C1(n8560), .C2(n9389), .A(n1755), 
        .ZN(n1748) );
  OAI221_X1 U807 ( .B1(n8496), .B2(n9404), .C1(n8257), .C2(n9401), .A(n1754), 
        .ZN(n1749) );
  OAI221_X1 U808 ( .B1(n8457), .B2(n9416), .C1(n8425), .C2(n9413), .A(n1753), 
        .ZN(n1750) );
  NOR4_X1 U809 ( .A1(n1730), .A2(n1731), .A3(n1732), .A4(n1733), .ZN(n1729) );
  OAI221_X1 U810 ( .B1(n8585), .B2(n9392), .C1(n8561), .C2(n9389), .A(n1737), 
        .ZN(n1730) );
  OAI221_X1 U811 ( .B1(n8497), .B2(n9404), .C1(n8258), .C2(n9401), .A(n1736), 
        .ZN(n1731) );
  OAI221_X1 U812 ( .B1(n8458), .B2(n9416), .C1(n8426), .C2(n9413), .A(n1735), 
        .ZN(n1732) );
  NOR4_X1 U813 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .ZN(n1711) );
  OAI221_X1 U814 ( .B1(n8586), .B2(n9392), .C1(n8562), .C2(n9389), .A(n1719), 
        .ZN(n1712) );
  OAI221_X1 U815 ( .B1(n8498), .B2(n9404), .C1(n8259), .C2(n9401), .A(n1718), 
        .ZN(n1713) );
  OAI221_X1 U816 ( .B1(n8459), .B2(n9416), .C1(n8427), .C2(n9413), .A(n1717), 
        .ZN(n1714) );
  NOR4_X1 U817 ( .A1(n1694), .A2(n1695), .A3(n1696), .A4(n1697), .ZN(n1693) );
  OAI221_X1 U818 ( .B1(n8587), .B2(n9392), .C1(n8563), .C2(n9389), .A(n1701), 
        .ZN(n1694) );
  OAI221_X1 U819 ( .B1(n8499), .B2(n9404), .C1(n8260), .C2(n9401), .A(n1700), 
        .ZN(n1695) );
  OAI221_X1 U820 ( .B1(n8460), .B2(n9416), .C1(n8428), .C2(n9413), .A(n1699), 
        .ZN(n1696) );
  NOR4_X1 U821 ( .A1(n1676), .A2(n1677), .A3(n1678), .A4(n1679), .ZN(n1675) );
  OAI221_X1 U822 ( .B1(n8588), .B2(n9392), .C1(n8564), .C2(n9389), .A(n1683), 
        .ZN(n1676) );
  OAI221_X1 U823 ( .B1(n8500), .B2(n9404), .C1(n8261), .C2(n9401), .A(n1682), 
        .ZN(n1677) );
  OAI221_X1 U824 ( .B1(n8461), .B2(n9416), .C1(n8429), .C2(n9413), .A(n1681), 
        .ZN(n1678) );
  NOR4_X1 U825 ( .A1(n1658), .A2(n1659), .A3(n1660), .A4(n1661), .ZN(n1657) );
  OAI221_X1 U826 ( .B1(n8589), .B2(n9392), .C1(n8565), .C2(n9389), .A(n1665), 
        .ZN(n1658) );
  OAI221_X1 U827 ( .B1(n8501), .B2(n9404), .C1(n8262), .C2(n9401), .A(n1664), 
        .ZN(n1659) );
  OAI221_X1 U828 ( .B1(n8462), .B2(n9416), .C1(n8430), .C2(n9413), .A(n1663), 
        .ZN(n1660) );
  NOR4_X1 U829 ( .A1(n1640), .A2(n1641), .A3(n1642), .A4(n1643), .ZN(n1639) );
  OAI221_X1 U830 ( .B1(n8590), .B2(n9393), .C1(n8319), .C2(n9390), .A(n1647), 
        .ZN(n1640) );
  OAI221_X1 U831 ( .B1(n8502), .B2(n9405), .C1(n8327), .C2(n9402), .A(n1646), 
        .ZN(n1641) );
  OAI221_X1 U832 ( .B1(n8463), .B2(n9417), .C1(n8431), .C2(n9414), .A(n1645), 
        .ZN(n1642) );
  NOR4_X1 U833 ( .A1(n1622), .A2(n1623), .A3(n1624), .A4(n1625), .ZN(n1621) );
  OAI221_X1 U834 ( .B1(n8591), .B2(n9393), .C1(n8320), .C2(n9390), .A(n1629), 
        .ZN(n1622) );
  OAI221_X1 U835 ( .B1(n8503), .B2(n9405), .C1(n8328), .C2(n9402), .A(n1628), 
        .ZN(n1623) );
  OAI221_X1 U836 ( .B1(n8464), .B2(n9417), .C1(n8432), .C2(n9414), .A(n1627), 
        .ZN(n1624) );
  NOR4_X1 U837 ( .A1(n1604), .A2(n1605), .A3(n1606), .A4(n1607), .ZN(n1603) );
  OAI221_X1 U838 ( .B1(n8592), .B2(n9393), .C1(n8321), .C2(n9390), .A(n1611), 
        .ZN(n1604) );
  OAI221_X1 U839 ( .B1(n8504), .B2(n9405), .C1(n8329), .C2(n9402), .A(n1610), 
        .ZN(n1605) );
  OAI221_X1 U840 ( .B1(n8465), .B2(n9417), .C1(n8433), .C2(n9414), .A(n1609), 
        .ZN(n1606) );
  NOR4_X1 U841 ( .A1(n1586), .A2(n1587), .A3(n1588), .A4(n1589), .ZN(n1585) );
  OAI221_X1 U842 ( .B1(n8593), .B2(n9393), .C1(n8322), .C2(n9390), .A(n1593), 
        .ZN(n1586) );
  OAI221_X1 U843 ( .B1(n8505), .B2(n9405), .C1(n8330), .C2(n9402), .A(n1592), 
        .ZN(n1587) );
  OAI221_X1 U844 ( .B1(n8466), .B2(n9417), .C1(n8434), .C2(n9414), .A(n1591), 
        .ZN(n1588) );
  NOR4_X1 U845 ( .A1(n1568), .A2(n1569), .A3(n1570), .A4(n1571), .ZN(n1567) );
  OAI221_X1 U846 ( .B1(n8594), .B2(n9393), .C1(n8323), .C2(n9390), .A(n1575), 
        .ZN(n1568) );
  OAI221_X1 U847 ( .B1(n8506), .B2(n9405), .C1(n8331), .C2(n9402), .A(n1574), 
        .ZN(n1569) );
  OAI221_X1 U848 ( .B1(n8467), .B2(n9417), .C1(n8435), .C2(n9414), .A(n1573), 
        .ZN(n1570) );
  NOR4_X1 U849 ( .A1(n1550), .A2(n1551), .A3(n1552), .A4(n1553), .ZN(n1549) );
  OAI221_X1 U850 ( .B1(n8595), .B2(n9393), .C1(n8324), .C2(n9390), .A(n1557), 
        .ZN(n1550) );
  OAI221_X1 U851 ( .B1(n8507), .B2(n9405), .C1(n8332), .C2(n9402), .A(n1556), 
        .ZN(n1551) );
  OAI221_X1 U852 ( .B1(n8468), .B2(n9417), .C1(n8436), .C2(n9414), .A(n1555), 
        .ZN(n1552) );
  NOR4_X1 U853 ( .A1(n1532), .A2(n1533), .A3(n1534), .A4(n1535), .ZN(n1531) );
  OAI221_X1 U854 ( .B1(n8596), .B2(n9393), .C1(n8325), .C2(n9390), .A(n1539), 
        .ZN(n1532) );
  OAI221_X1 U855 ( .B1(n8508), .B2(n9405), .C1(n8333), .C2(n9402), .A(n1538), 
        .ZN(n1533) );
  OAI221_X1 U856 ( .B1(n8469), .B2(n9417), .C1(n8437), .C2(n9414), .A(n1537), 
        .ZN(n1534) );
  NOR4_X1 U857 ( .A1(n1482), .A2(n1483), .A3(n1484), .A4(n1485), .ZN(n1481) );
  OAI221_X1 U858 ( .B1(n8597), .B2(n9393), .C1(n8326), .C2(n9390), .A(n1503), 
        .ZN(n1482) );
  OAI221_X1 U859 ( .B1(n8509), .B2(n9405), .C1(n8334), .C2(n9402), .A(n1498), 
        .ZN(n1483) );
  OAI221_X1 U860 ( .B1(n8470), .B2(n9417), .C1(n8438), .C2(n9414), .A(n1493), 
        .ZN(n1484) );
  NOR4_X1 U861 ( .A1(n2090), .A2(n2091), .A3(n2092), .A4(n2093), .ZN(n2070) );
  OAI221_X1 U862 ( .B1(n8886), .B2(n9343), .C1(n8862), .C2(n9340), .A(n2099), 
        .ZN(n2090) );
  OAI221_X1 U863 ( .B1(n8742), .B2(n9367), .C1(n8718), .C2(n9364), .A(n2096), 
        .ZN(n2092) );
  OAI221_X1 U864 ( .B1(n8798), .B2(n9355), .C1(n8774), .C2(n9352), .A(n2097), 
        .ZN(n2091) );
  NOR4_X1 U865 ( .A1(n2062), .A2(n2063), .A3(n2064), .A4(n2065), .ZN(n2052) );
  OAI221_X1 U866 ( .B1(n8887), .B2(n9343), .C1(n8863), .C2(n9340), .A(n2069), 
        .ZN(n2062) );
  OAI221_X1 U867 ( .B1(n8743), .B2(n9367), .C1(n8719), .C2(n9364), .A(n2067), 
        .ZN(n2064) );
  OAI221_X1 U868 ( .B1(n8799), .B2(n9355), .C1(n8775), .C2(n9352), .A(n2068), 
        .ZN(n2063) );
  NOR4_X1 U869 ( .A1(n2044), .A2(n2045), .A3(n2046), .A4(n2047), .ZN(n2034) );
  OAI221_X1 U870 ( .B1(n8888), .B2(n9343), .C1(n8864), .C2(n9340), .A(n2051), 
        .ZN(n2044) );
  OAI221_X1 U871 ( .B1(n8744), .B2(n9367), .C1(n8720), .C2(n9364), .A(n2049), 
        .ZN(n2046) );
  OAI221_X1 U872 ( .B1(n8800), .B2(n9355), .C1(n8776), .C2(n9352), .A(n2050), 
        .ZN(n2045) );
  NOR4_X1 U873 ( .A1(n2026), .A2(n2027), .A3(n2028), .A4(n2029), .ZN(n2016) );
  OAI221_X1 U874 ( .B1(n8889), .B2(n9343), .C1(n8865), .C2(n9340), .A(n2033), 
        .ZN(n2026) );
  OAI221_X1 U875 ( .B1(n8745), .B2(n9367), .C1(n8721), .C2(n9364), .A(n2031), 
        .ZN(n2028) );
  OAI221_X1 U876 ( .B1(n8801), .B2(n9355), .C1(n8777), .C2(n9352), .A(n2032), 
        .ZN(n2027) );
  NOR4_X1 U877 ( .A1(n2008), .A2(n2009), .A3(n2010), .A4(n2011), .ZN(n1998) );
  OAI221_X1 U878 ( .B1(n8890), .B2(n9343), .C1(n8866), .C2(n9340), .A(n2015), 
        .ZN(n2008) );
  OAI221_X1 U879 ( .B1(n8746), .B2(n9367), .C1(n8722), .C2(n9364), .A(n2013), 
        .ZN(n2010) );
  OAI221_X1 U880 ( .B1(n8802), .B2(n9355), .C1(n8778), .C2(n9352), .A(n2014), 
        .ZN(n2009) );
  NOR4_X1 U881 ( .A1(n1990), .A2(n1991), .A3(n1992), .A4(n1993), .ZN(n1980) );
  OAI221_X1 U882 ( .B1(n8891), .B2(n9343), .C1(n8867), .C2(n9340), .A(n1997), 
        .ZN(n1990) );
  OAI221_X1 U883 ( .B1(n8747), .B2(n9367), .C1(n8723), .C2(n9364), .A(n1995), 
        .ZN(n1992) );
  OAI221_X1 U884 ( .B1(n8803), .B2(n9355), .C1(n8779), .C2(n9352), .A(n1996), 
        .ZN(n1991) );
  NOR4_X1 U885 ( .A1(n1972), .A2(n1973), .A3(n1974), .A4(n1975), .ZN(n1962) );
  OAI221_X1 U886 ( .B1(n8892), .B2(n9343), .C1(n8868), .C2(n9340), .A(n1979), 
        .ZN(n1972) );
  OAI221_X1 U887 ( .B1(n8748), .B2(n9367), .C1(n8724), .C2(n9364), .A(n1977), 
        .ZN(n1974) );
  OAI221_X1 U888 ( .B1(n8804), .B2(n9355), .C1(n8780), .C2(n9352), .A(n1978), 
        .ZN(n1973) );
  NOR4_X1 U889 ( .A1(n1954), .A2(n1955), .A3(n1956), .A4(n1957), .ZN(n1944) );
  OAI221_X1 U890 ( .B1(n8893), .B2(n9343), .C1(n8869), .C2(n9340), .A(n1961), 
        .ZN(n1954) );
  OAI221_X1 U891 ( .B1(n8749), .B2(n9367), .C1(n8725), .C2(n9364), .A(n1959), 
        .ZN(n1956) );
  OAI221_X1 U892 ( .B1(n8805), .B2(n9355), .C1(n8781), .C2(n9352), .A(n1960), 
        .ZN(n1955) );
  NAND2_X1 U893 ( .A1(n982), .A2(n983), .ZN(N716) );
  NOR4_X1 U894 ( .A1(n984), .A2(n985), .A3(n986), .A4(n987), .ZN(n983) );
  NOR4_X1 U895 ( .A1(n992), .A2(n993), .A3(n994), .A4(n995), .ZN(n982) );
  OAI221_X1 U896 ( .B1(n2143), .B2(n9489), .C1(n8401), .C2(n9486), .A(n991), 
        .ZN(n984) );
  AND3_X1 U897 ( .A1(n849), .A2(n9918), .A3(ADD_WR[4]), .ZN(n816) );
  AND3_X1 U898 ( .A1(ADD_WR[4]), .A2(n849), .A3(ADD_WR[3]), .ZN(n821) );
  AND3_X1 U899 ( .A1(n849), .A2(n9917), .A3(ADD_WR[3]), .ZN(n826) );
  OAI221_X1 U900 ( .B1(n8658), .B2(n9475), .C1(n8634), .C2(n9472), .A(n1392), 
        .ZN(n1391) );
  AOI22_X1 U901 ( .A1(n9469), .A2(n10189), .B1(n9468), .B2(n10253), .ZN(n1392)
         );
  OAI221_X1 U902 ( .B1(n8659), .B2(n9475), .C1(n8635), .C2(n9472), .A(n1374), 
        .ZN(n1373) );
  AOI22_X1 U903 ( .A1(n9469), .A2(n10188), .B1(n9468), .B2(n10252), .ZN(n1374)
         );
  OAI221_X1 U904 ( .B1(n8674), .B2(n9476), .C1(n8650), .C2(n9473), .A(n1104), 
        .ZN(n1103) );
  AOI22_X1 U905 ( .A1(n9470), .A2(n10173), .B1(n9466), .B2(n10237), .ZN(n1104)
         );
  OAI221_X1 U906 ( .B1(n8669), .B2(n9476), .C1(n8645), .C2(n9473), .A(n1194), 
        .ZN(n1193) );
  AOI22_X1 U907 ( .A1(n9470), .A2(n10178), .B1(n9467), .B2(n10242), .ZN(n1194)
         );
  OAI221_X1 U908 ( .B1(n8675), .B2(n9476), .C1(n8651), .C2(n9473), .A(n1086), 
        .ZN(n1085) );
  AOI22_X1 U909 ( .A1(n9470), .A2(n10172), .B1(n9466), .B2(n10236), .ZN(n1086)
         );
  OAI221_X1 U910 ( .B1(n8665), .B2(n9475), .C1(n8641), .C2(n9472), .A(n1266), 
        .ZN(n1265) );
  AOI22_X1 U911 ( .A1(n9469), .A2(n10182), .B1(n9467), .B2(n10246), .ZN(n1266)
         );
  OAI221_X1 U912 ( .B1(n8676), .B2(n9476), .C1(n8652), .C2(n9473), .A(n1068), 
        .ZN(n1067) );
  AOI22_X1 U913 ( .A1(n9470), .A2(n10171), .B1(n9466), .B2(n10235), .ZN(n1068)
         );
  OAI221_X1 U914 ( .B1(n8670), .B2(n9476), .C1(n8646), .C2(n9473), .A(n1176), 
        .ZN(n1175) );
  AOI22_X1 U915 ( .A1(n9470), .A2(n10177), .B1(n9467), .B2(n10241), .ZN(n1176)
         );
  OAI221_X1 U916 ( .B1(n8666), .B2(n9476), .C1(n8642), .C2(n9473), .A(n1248), 
        .ZN(n1247) );
  AOI22_X1 U917 ( .A1(n9470), .A2(n10181), .B1(n9467), .B2(n10245), .ZN(n1248)
         );
  OAI221_X1 U918 ( .B1(n8677), .B2(n9476), .C1(n8653), .C2(n9473), .A(n1050), 
        .ZN(n1049) );
  AOI22_X1 U919 ( .A1(n9470), .A2(n10170), .B1(n9466), .B2(n10234), .ZN(n1050)
         );
  OAI221_X1 U920 ( .B1(n8673), .B2(n9476), .C1(n8649), .C2(n9473), .A(n1122), 
        .ZN(n1121) );
  AOI22_X1 U921 ( .A1(n9470), .A2(n10174), .B1(n9467), .B2(n10238), .ZN(n1122)
         );
  OAI221_X1 U922 ( .B1(n8655), .B2(n9475), .C1(n8631), .C2(n9472), .A(n1446), 
        .ZN(n1445) );
  AOI22_X1 U923 ( .A1(n9469), .A2(n10192), .B1(n9468), .B2(n10256), .ZN(n1446)
         );
  OAI221_X1 U924 ( .B1(n8679), .B2(n9477), .C1(n8296), .C2(n9474), .A(n1014), 
        .ZN(n1013) );
  AOI22_X1 U925 ( .A1(n9471), .A2(n10584), .B1(n9466), .B2(n10232), .ZN(n1014)
         );
  OAI221_X1 U926 ( .B1(n8656), .B2(n9475), .C1(n8632), .C2(n9472), .A(n1428), 
        .ZN(n1427) );
  AOI22_X1 U927 ( .A1(n9469), .A2(n10191), .B1(n9468), .B2(n10255), .ZN(n1428)
         );
  OAI221_X1 U928 ( .B1(n8661), .B2(n9475), .C1(n8637), .C2(n9472), .A(n1338), 
        .ZN(n1337) );
  AOI22_X1 U929 ( .A1(n9469), .A2(n10186), .B1(n9468), .B2(n10250), .ZN(n1338)
         );
  OAI221_X1 U930 ( .B1(n8680), .B2(n9477), .C1(n8297), .C2(n9474), .A(n996), 
        .ZN(n995) );
  AOI22_X1 U931 ( .A1(n9471), .A2(n10583), .B1(n9466), .B2(n10231), .ZN(n996)
         );
  OAI221_X1 U932 ( .B1(n8662), .B2(n9475), .C1(n8638), .C2(n9472), .A(n1320), 
        .ZN(n1319) );
  AOI22_X1 U933 ( .A1(n9469), .A2(n10185), .B1(n9467), .B2(n10249), .ZN(n1320)
         );
  OAI221_X1 U934 ( .B1(n8684), .B2(n9477), .C1(n8301), .C2(n9474), .A(n924), 
        .ZN(n923) );
  AOI22_X1 U935 ( .A1(n9471), .A2(n10579), .B1(n9466), .B2(n10227), .ZN(n924)
         );
  OAI221_X1 U936 ( .B1(n8681), .B2(n9477), .C1(n8298), .C2(n9474), .A(n978), 
        .ZN(n977) );
  AOI22_X1 U937 ( .A1(n9471), .A2(n10582), .B1(n9466), .B2(n10230), .ZN(n978)
         );
  OAI221_X1 U938 ( .B1(n8663), .B2(n9475), .C1(n8639), .C2(n9472), .A(n1302), 
        .ZN(n1301) );
  AOI22_X1 U939 ( .A1(n9469), .A2(n10184), .B1(n9467), .B2(n10248), .ZN(n1302)
         );
  OAI221_X1 U940 ( .B1(n8662), .B2(n9379), .C1(n8638), .C2(n9376), .A(n1940), 
        .ZN(n1939) );
  AOI22_X1 U941 ( .A1(n9373), .A2(n10217), .B1(n9371), .B2(n10249), .ZN(n1940)
         );
  OAI221_X1 U942 ( .B1(n8663), .B2(n9379), .C1(n8639), .C2(n9376), .A(n1922), 
        .ZN(n1921) );
  AOI22_X1 U943 ( .A1(n9373), .A2(n10216), .B1(n9371), .B2(n10248), .ZN(n1922)
         );
  OAI221_X1 U944 ( .B1(n8664), .B2(n9379), .C1(n8640), .C2(n9376), .A(n1904), 
        .ZN(n1903) );
  AOI22_X1 U945 ( .A1(n9373), .A2(n10215), .B1(n9371), .B2(n10247), .ZN(n1904)
         );
  OAI221_X1 U946 ( .B1(n8665), .B2(n9379), .C1(n8641), .C2(n9376), .A(n1886), 
        .ZN(n1885) );
  AOI22_X1 U947 ( .A1(n9373), .A2(n10214), .B1(n9371), .B2(n10246), .ZN(n1886)
         );
  OAI221_X1 U948 ( .B1(n8666), .B2(n9380), .C1(n8642), .C2(n9377), .A(n1868), 
        .ZN(n1867) );
  AOI22_X1 U949 ( .A1(n9374), .A2(n10213), .B1(n9371), .B2(n10245), .ZN(n1868)
         );
  OAI221_X1 U950 ( .B1(n8668), .B2(n9380), .C1(n8644), .C2(n9377), .A(n1832), 
        .ZN(n1831) );
  AOI22_X1 U951 ( .A1(n9374), .A2(n10211), .B1(n9371), .B2(n10243), .ZN(n1832)
         );
  OAI221_X1 U952 ( .B1(n8669), .B2(n9380), .C1(n8645), .C2(n9377), .A(n1814), 
        .ZN(n1813) );
  AOI22_X1 U953 ( .A1(n9374), .A2(n10210), .B1(n9371), .B2(n10242), .ZN(n1814)
         );
  OAI221_X1 U954 ( .B1(n8670), .B2(n9380), .C1(n8646), .C2(n9377), .A(n1796), 
        .ZN(n1795) );
  AOI22_X1 U955 ( .A1(n9374), .A2(n10209), .B1(n9371), .B2(n10241), .ZN(n1796)
         );
  OAI221_X1 U956 ( .B1(n8672), .B2(n9380), .C1(n8648), .C2(n9377), .A(n1760), 
        .ZN(n1759) );
  AOI22_X1 U957 ( .A1(n9374), .A2(n10207), .B1(n9371), .B2(n10239), .ZN(n1760)
         );
  OAI221_X1 U958 ( .B1(n8673), .B2(n9380), .C1(n8649), .C2(n9377), .A(n1742), 
        .ZN(n1741) );
  AOI22_X1 U959 ( .A1(n9374), .A2(n10206), .B1(n9371), .B2(n10238), .ZN(n1742)
         );
  OAI221_X1 U960 ( .B1(n8674), .B2(n9380), .C1(n8650), .C2(n9377), .A(n1724), 
        .ZN(n1723) );
  AOI22_X1 U961 ( .A1(n9374), .A2(n10205), .B1(n9370), .B2(n10237), .ZN(n1724)
         );
  OAI221_X1 U962 ( .B1(n8675), .B2(n9380), .C1(n8651), .C2(n9377), .A(n1706), 
        .ZN(n1705) );
  AOI22_X1 U963 ( .A1(n9374), .A2(n10204), .B1(n9370), .B2(n10236), .ZN(n1706)
         );
  OAI221_X1 U964 ( .B1(n8676), .B2(n9380), .C1(n8652), .C2(n9377), .A(n1688), 
        .ZN(n1687) );
  AOI22_X1 U965 ( .A1(n9374), .A2(n10203), .B1(n9370), .B2(n10235), .ZN(n1688)
         );
  OAI221_X1 U966 ( .B1(n8677), .B2(n9380), .C1(n8653), .C2(n9377), .A(n1670), 
        .ZN(n1669) );
  AOI22_X1 U967 ( .A1(n9374), .A2(n10202), .B1(n9370), .B2(n10234), .ZN(n1670)
         );
  OAI221_X1 U968 ( .B1(n8678), .B2(n9381), .C1(n8295), .C2(n9378), .A(n1652), 
        .ZN(n1651) );
  AOI22_X1 U969 ( .A1(n9375), .A2(n10201), .B1(n9370), .B2(n10233), .ZN(n1652)
         );
  OAI221_X1 U970 ( .B1(n8679), .B2(n9381), .C1(n8296), .C2(n9378), .A(n1634), 
        .ZN(n1633) );
  AOI22_X1 U971 ( .A1(n9375), .A2(n10200), .B1(n9370), .B2(n10232), .ZN(n1634)
         );
  OAI221_X1 U972 ( .B1(n8680), .B2(n9381), .C1(n8297), .C2(n9378), .A(n1616), 
        .ZN(n1615) );
  AOI22_X1 U973 ( .A1(n9375), .A2(n10199), .B1(n9370), .B2(n10231), .ZN(n1616)
         );
  OAI221_X1 U974 ( .B1(n8681), .B2(n9381), .C1(n8298), .C2(n9378), .A(n1598), 
        .ZN(n1597) );
  AOI22_X1 U975 ( .A1(n9375), .A2(n10198), .B1(n9370), .B2(n10230), .ZN(n1598)
         );
  OAI221_X1 U976 ( .B1(n8682), .B2(n9381), .C1(n8299), .C2(n9378), .A(n1580), 
        .ZN(n1579) );
  AOI22_X1 U977 ( .A1(n9375), .A2(n10197), .B1(n9370), .B2(n10229), .ZN(n1580)
         );
  OAI221_X1 U978 ( .B1(n8683), .B2(n9381), .C1(n8300), .C2(n9378), .A(n1562), 
        .ZN(n1561) );
  AOI22_X1 U979 ( .A1(n9375), .A2(n10196), .B1(n9370), .B2(n10228), .ZN(n1562)
         );
  OAI221_X1 U980 ( .B1(n8684), .B2(n9381), .C1(n8301), .C2(n9378), .A(n1544), 
        .ZN(n1543) );
  AOI22_X1 U981 ( .A1(n9375), .A2(n10195), .B1(n9370), .B2(n10227), .ZN(n1544)
         );
  OAI221_X1 U982 ( .B1(n8685), .B2(n9381), .C1(n8302), .C2(n9378), .A(n1512), 
        .ZN(n1509) );
  AOI22_X1 U983 ( .A1(n9375), .A2(n10194), .B1(n9370), .B2(n10226), .ZN(n1512)
         );
  OAI221_X1 U984 ( .B1(n8601), .B2(n9523), .C1(n8569), .C2(n9520), .A(n1402), 
        .ZN(n1401) );
  AOI22_X1 U985 ( .A1(n9517), .A2(n10470), .B1(n9516), .B2(n10286), .ZN(n1402)
         );
  OAI221_X1 U986 ( .B1(n8602), .B2(n9523), .C1(n8570), .C2(n9520), .A(n1384), 
        .ZN(n1383) );
  AOI22_X1 U987 ( .A1(n9517), .A2(n10469), .B1(n9516), .B2(n10285), .ZN(n1384)
         );
  OAI221_X1 U988 ( .B1(n8603), .B2(n9523), .C1(n8571), .C2(n9520), .A(n1366), 
        .ZN(n1365) );
  AOI22_X1 U989 ( .A1(n9517), .A2(n10468), .B1(n9516), .B2(n10284), .ZN(n1366)
         );
  OAI221_X1 U990 ( .B1(n8618), .B2(n9524), .C1(n8586), .C2(n9521), .A(n1096), 
        .ZN(n1095) );
  AOI22_X1 U991 ( .A1(n9518), .A2(n10453), .B1(n9514), .B2(n10269), .ZN(n1096)
         );
  OAI221_X1 U992 ( .B1(n8608), .B2(n9523), .C1(n8576), .C2(n9520), .A(n1276), 
        .ZN(n1275) );
  AOI22_X1 U993 ( .A1(n9517), .A2(n10463), .B1(n9515), .B2(n10279), .ZN(n1276)
         );
  OAI221_X1 U994 ( .B1(n8609), .B2(n9523), .C1(n8577), .C2(n9520), .A(n1258), 
        .ZN(n1257) );
  AOI22_X1 U995 ( .A1(n9517), .A2(n10462), .B1(n9515), .B2(n10278), .ZN(n1258)
         );
  OAI221_X1 U996 ( .B1(n8620), .B2(n9524), .C1(n8588), .C2(n9521), .A(n1060), 
        .ZN(n1059) );
  AOI22_X1 U997 ( .A1(n9518), .A2(n10451), .B1(n9514), .B2(n10267), .ZN(n1060)
         );
  OAI221_X1 U998 ( .B1(n8619), .B2(n9524), .C1(n8587), .C2(n9521), .A(n1078), 
        .ZN(n1077) );
  AOI22_X1 U999 ( .A1(n9518), .A2(n10452), .B1(n9514), .B2(n10268), .ZN(n1078)
         );
  OAI221_X1 U1000 ( .B1(n8614), .B2(n9524), .C1(n8582), .C2(n9521), .A(n1168), 
        .ZN(n1167) );
  AOI22_X1 U1001 ( .A1(n9518), .A2(n10457), .B1(n9515), .B2(n10273), .ZN(n1168) );
  OAI221_X1 U1002 ( .B1(n8610), .B2(n9524), .C1(n8578), .C2(n9521), .A(n1240), 
        .ZN(n1239) );
  AOI22_X1 U1003 ( .A1(n9518), .A2(n10461), .B1(n9515), .B2(n10277), .ZN(n1240) );
  OAI221_X1 U1004 ( .B1(n8621), .B2(n9524), .C1(n8589), .C2(n9521), .A(n1042), 
        .ZN(n1041) );
  AOI22_X1 U1005 ( .A1(n9518), .A2(n10450), .B1(n9514), .B2(n10266), .ZN(n1042) );
  OAI221_X1 U1006 ( .B1(n8599), .B2(n9523), .C1(n8567), .C2(n9520), .A(n1438), 
        .ZN(n1437) );
  AOI22_X1 U1007 ( .A1(n9517), .A2(n10472), .B1(n9516), .B2(n10288), .ZN(n1438) );
  OAI221_X1 U1008 ( .B1(n8600), .B2(n9523), .C1(n8568), .C2(n9520), .A(n1420), 
        .ZN(n1419) );
  AOI22_X1 U1009 ( .A1(n9517), .A2(n10471), .B1(n9516), .B2(n10287), .ZN(n1420) );
  OAI221_X1 U1010 ( .B1(n8604), .B2(n9523), .C1(n8572), .C2(n9520), .A(n1348), 
        .ZN(n1347) );
  AOI22_X1 U1011 ( .A1(n9517), .A2(n10467), .B1(n9516), .B2(n10283), .ZN(n1348) );
  OAI221_X1 U1012 ( .B1(n8622), .B2(n9525), .C1(n8590), .C2(n9522), .A(n1024), 
        .ZN(n1023) );
  AOI22_X1 U1013 ( .A1(n9519), .A2(n10449), .B1(n9514), .B2(n10265), .ZN(n1024) );
  OAI221_X1 U1014 ( .B1(n8627), .B2(n9525), .C1(n8595), .C2(n9522), .A(n934), 
        .ZN(n933) );
  AOI22_X1 U1015 ( .A1(n9519), .A2(n10444), .B1(n9514), .B2(n10260), .ZN(n934)
         );
  OAI221_X1 U1016 ( .B1(n8605), .B2(n9523), .C1(n8573), .C2(n9520), .A(n1330), 
        .ZN(n1329) );
  AOI22_X1 U1017 ( .A1(n9517), .A2(n10466), .B1(n9516), .B2(n10282), .ZN(n1330) );
  OAI221_X1 U1018 ( .B1(n8624), .B2(n9525), .C1(n8592), .C2(n9522), .A(n988), 
        .ZN(n987) );
  AOI22_X1 U1019 ( .A1(n9519), .A2(n10447), .B1(n9514), .B2(n10263), .ZN(n988)
         );
  OAI221_X1 U1020 ( .B1(n8628), .B2(n9525), .C1(n8596), .C2(n9522), .A(n916), 
        .ZN(n915) );
  AOI22_X1 U1021 ( .A1(n9519), .A2(n10443), .B1(n9514), .B2(n10259), .ZN(n916)
         );
  OAI221_X1 U1022 ( .B1(n8606), .B2(n9523), .C1(n8574), .C2(n9520), .A(n1312), 
        .ZN(n1311) );
  AOI22_X1 U1023 ( .A1(n9517), .A2(n10465), .B1(n9515), .B2(n10281), .ZN(n1312) );
  OAI221_X1 U1024 ( .B1(n8625), .B2(n9525), .C1(n8593), .C2(n9522), .A(n970), 
        .ZN(n969) );
  AOI22_X1 U1025 ( .A1(n9519), .A2(n10446), .B1(n9514), .B2(n10262), .ZN(n970)
         );
  OAI221_X1 U1026 ( .B1(n8607), .B2(n9523), .C1(n8575), .C2(n9520), .A(n1294), 
        .ZN(n1293) );
  AOI22_X1 U1027 ( .A1(n9517), .A2(n10464), .B1(n9515), .B2(n10280), .ZN(n1294) );
  OAI221_X1 U1028 ( .B1(n8667), .B2(n9380), .C1(n8643), .C2(n9377), .A(n1850), 
        .ZN(n1849) );
  AOI22_X1 U1029 ( .A1(n9374), .A2(n10212), .B1(n9371), .B2(n10244), .ZN(n1850) );
  OAI221_X1 U1030 ( .B1(n8671), .B2(n9380), .C1(n8647), .C2(n9377), .A(n1778), 
        .ZN(n1777) );
  AOI22_X1 U1031 ( .A1(n9374), .A2(n10208), .B1(n9371), .B2(n10240), .ZN(n1778) );
  OAI221_X1 U1032 ( .B1(n8778), .B2(n9463), .C1(n8237), .C2(n9460), .A(n1393), 
        .ZN(n1390) );
  AOI22_X1 U1033 ( .A1(n9457), .A2(n10133), .B1(n9456), .B2(n10165), .ZN(n1393) );
  OAI221_X1 U1034 ( .B1(n8334), .B2(n9513), .C1(n8182), .C2(n9510), .A(n873), 
        .ZN(n864) );
  AOI22_X1 U1035 ( .A1(n9507), .A2(n10538), .B1(n9502), .B2(n10410), .ZN(n873)
         );
  OAI221_X1 U1036 ( .B1(n8779), .B2(n9463), .C1(n8235), .C2(n9460), .A(n1375), 
        .ZN(n1372) );
  AOI22_X1 U1037 ( .A1(n9457), .A2(n10132), .B1(n9456), .B2(n10164), .ZN(n1375) );
  OAI221_X1 U1038 ( .B1(n8794), .B2(n9464), .C1(n8205), .C2(n9461), .A(n1105), 
        .ZN(n1102) );
  AOI22_X1 U1039 ( .A1(n9458), .A2(n10117), .B1(n9454), .B2(n10149), .ZN(n1105) );
  OAI221_X1 U1040 ( .B1(n8789), .B2(n9464), .C1(n8215), .C2(n9461), .A(n1195), 
        .ZN(n1192) );
  AOI22_X1 U1041 ( .A1(n9458), .A2(n10122), .B1(n9455), .B2(n10154), .ZN(n1195) );
  OAI221_X1 U1042 ( .B1(n8795), .B2(n9464), .C1(n8203), .C2(n9461), .A(n1087), 
        .ZN(n1084) );
  AOI22_X1 U1043 ( .A1(n9458), .A2(n10116), .B1(n9454), .B2(n10148), .ZN(n1087) );
  OAI221_X1 U1044 ( .B1(n8785), .B2(n9463), .C1(n8223), .C2(n9460), .A(n1267), 
        .ZN(n1264) );
  AOI22_X1 U1045 ( .A1(n9457), .A2(n10126), .B1(n9455), .B2(n10158), .ZN(n1267) );
  OAI221_X1 U1046 ( .B1(n8796), .B2(n9464), .C1(n8201), .C2(n9461), .A(n1069), 
        .ZN(n1066) );
  AOI22_X1 U1047 ( .A1(n9458), .A2(n10115), .B1(n9454), .B2(n10147), .ZN(n1069) );
  OAI221_X1 U1048 ( .B1(n8471), .B2(n9511), .C1(n8244), .C2(n9508), .A(n1462), 
        .ZN(n1454) );
  AOI22_X1 U1049 ( .A1(n9505), .A2(n10609), .B1(n9504), .B2(n10441), .ZN(n1462) );
  OAI221_X1 U1050 ( .B1(n8790), .B2(n9464), .C1(n8213), .C2(n9461), .A(n1177), 
        .ZN(n1174) );
  AOI22_X1 U1051 ( .A1(n9458), .A2(n10121), .B1(n9455), .B2(n10153), .ZN(n1177) );
  OAI221_X1 U1052 ( .B1(n8786), .B2(n9464), .C1(n8221), .C2(n9461), .A(n1249), 
        .ZN(n1246) );
  AOI22_X1 U1053 ( .A1(n9458), .A2(n10125), .B1(n9455), .B2(n10157), .ZN(n1249) );
  OAI221_X1 U1054 ( .B1(n8797), .B2(n9464), .C1(n8199), .C2(n9461), .A(n1051), 
        .ZN(n1048) );
  AOI22_X1 U1055 ( .A1(n9458), .A2(n10114), .B1(n9454), .B2(n10146), .ZN(n1051) );
  OAI221_X1 U1056 ( .B1(n8793), .B2(n9464), .C1(n8207), .C2(n9461), .A(n1123), 
        .ZN(n1120) );
  AOI22_X1 U1057 ( .A1(n9458), .A2(n10118), .B1(n9455), .B2(n10150), .ZN(n1123) );
  OAI221_X1 U1058 ( .B1(n8775), .B2(n9463), .C1(n8243), .C2(n9460), .A(n1447), 
        .ZN(n1444) );
  AOI22_X1 U1059 ( .A1(n9457), .A2(n10136), .B1(n9456), .B2(n10168), .ZN(n1447) );
  OAI221_X1 U1060 ( .B1(n8312), .B2(n9465), .C1(n8195), .C2(n9462), .A(n1015), 
        .ZN(n1012) );
  AOI22_X1 U1061 ( .A1(n9459), .A2(n10112), .B1(n9454), .B2(n10144), .ZN(n1015) );
  OAI221_X1 U1062 ( .B1(n8776), .B2(n9463), .C1(n8241), .C2(n9460), .A(n1429), 
        .ZN(n1426) );
  AOI22_X1 U1063 ( .A1(n9457), .A2(n10135), .B1(n9456), .B2(n10167), .ZN(n1429) );
  OAI221_X1 U1064 ( .B1(n8781), .B2(n9463), .C1(n8231), .C2(n9460), .A(n1339), 
        .ZN(n1336) );
  AOI22_X1 U1065 ( .A1(n9457), .A2(n10130), .B1(n9456), .B2(n10162), .ZN(n1339) );
  OAI221_X1 U1066 ( .B1(n8313), .B2(n9465), .C1(n8193), .C2(n9462), .A(n997), 
        .ZN(n994) );
  AOI22_X1 U1067 ( .A1(n9459), .A2(n10111), .B1(n9454), .B2(n10143), .ZN(n997)
         );
  OAI221_X1 U1068 ( .B1(n8328), .B2(n9513), .C1(n8194), .C2(n9510), .A(n1007), 
        .ZN(n1004) );
  AOI22_X1 U1069 ( .A1(n9507), .A2(n10544), .B1(n9502), .B2(n10416), .ZN(n1007) );
  OAI221_X1 U1070 ( .B1(n8331), .B2(n9513), .C1(n8188), .C2(n9510), .A(n953), 
        .ZN(n950) );
  AOI22_X1 U1071 ( .A1(n9507), .A2(n10541), .B1(n9502), .B2(n10413), .ZN(n953)
         );
  OAI221_X1 U1072 ( .B1(n8327), .B2(n9513), .C1(n8196), .C2(n9510), .A(n1025), 
        .ZN(n1022) );
  AOI22_X1 U1073 ( .A1(n9507), .A2(n10545), .B1(n9502), .B2(n10417), .ZN(n1025) );
  OAI221_X1 U1074 ( .B1(n8332), .B2(n9513), .C1(n8186), .C2(n9510), .A(n935), 
        .ZN(n932) );
  AOI22_X1 U1075 ( .A1(n9507), .A2(n10540), .B1(n9502), .B2(n10412), .ZN(n935)
         );
  OAI221_X1 U1076 ( .B1(n8782), .B2(n9463), .C1(n8229), .C2(n9460), .A(n1321), 
        .ZN(n1318) );
  AOI22_X1 U1077 ( .A1(n9457), .A2(n10129), .B1(n9455), .B2(n10161), .ZN(n1321) );
  OAI221_X1 U1078 ( .B1(n8317), .B2(n9465), .C1(n8185), .C2(n9462), .A(n925), 
        .ZN(n922) );
  AOI22_X1 U1079 ( .A1(n9459), .A2(n10107), .B1(n9454), .B2(n10139), .ZN(n925)
         );
  OAI221_X1 U1080 ( .B1(n8329), .B2(n9513), .C1(n8192), .C2(n9510), .A(n989), 
        .ZN(n986) );
  AOI22_X1 U1081 ( .A1(n9507), .A2(n10543), .B1(n9502), .B2(n10415), .ZN(n989)
         );
  OAI221_X1 U1082 ( .B1(n8314), .B2(n9465), .C1(n8191), .C2(n9462), .A(n979), 
        .ZN(n976) );
  AOI22_X1 U1083 ( .A1(n9459), .A2(n10110), .B1(n9454), .B2(n10142), .ZN(n979)
         );
  OAI221_X1 U1084 ( .B1(n8783), .B2(n9463), .C1(n8227), .C2(n9460), .A(n1303), 
        .ZN(n1300) );
  AOI22_X1 U1085 ( .A1(n9457), .A2(n10128), .B1(n9455), .B2(n10160), .ZN(n1303) );
  OAI221_X1 U1086 ( .B1(n8477), .B2(n9511), .C1(n8232), .C2(n9508), .A(n1349), 
        .ZN(n1346) );
  AOI22_X1 U1087 ( .A1(n9505), .A2(n10603), .B1(n9504), .B2(n10435), .ZN(n1349) );
  OAI221_X1 U1088 ( .B1(n8333), .B2(n9513), .C1(n8184), .C2(n9510), .A(n917), 
        .ZN(n914) );
  AOI22_X1 U1089 ( .A1(n9507), .A2(n10539), .B1(n9502), .B2(n10411), .ZN(n917)
         );
  OAI221_X1 U1090 ( .B1(n8330), .B2(n9513), .C1(n8190), .C2(n9510), .A(n971), 
        .ZN(n968) );
  AOI22_X1 U1091 ( .A1(n9507), .A2(n10542), .B1(n9502), .B2(n10414), .ZN(n971)
         );
  OAI221_X1 U1092 ( .B1(n8513), .B2(n9499), .C1(n8481), .C2(n9496), .A(n1404), 
        .ZN(n1399) );
  AOI22_X1 U1093 ( .A1(n9493), .A2(n10502), .B1(n9492), .B2(n10374), .ZN(n1404) );
  OAI221_X1 U1094 ( .B1(n8541), .B2(n9501), .C1(n8509), .C2(n9498), .A(n878), 
        .ZN(n863) );
  AOI22_X1 U1095 ( .A1(n9495), .A2(n10474), .B1(n9490), .B2(n10346), .ZN(n878)
         );
  OAI221_X1 U1096 ( .B1(n8514), .B2(n9499), .C1(n8482), .C2(n9496), .A(n1386), 
        .ZN(n1381) );
  AOI22_X1 U1097 ( .A1(n9493), .A2(n10501), .B1(n9492), .B2(n10373), .ZN(n1386) );
  OAI221_X1 U1098 ( .B1(n8834), .B2(n9451), .C1(n8802), .C2(n9448), .A(n1394), 
        .ZN(n1389) );
  AOI22_X1 U1099 ( .A1(n9445), .A2(n10005), .B1(n9444), .B2(n10037), .ZN(n1394) );
  OAI221_X1 U1100 ( .B1(n8515), .B2(n9499), .C1(n8483), .C2(n9496), .A(n1368), 
        .ZN(n1363) );
  AOI22_X1 U1101 ( .A1(n9493), .A2(n10500), .B1(n9492), .B2(n10372), .ZN(n1368) );
  OAI221_X1 U1102 ( .B1(n8835), .B2(n9451), .C1(n8803), .C2(n9448), .A(n1376), 
        .ZN(n1371) );
  AOI22_X1 U1103 ( .A1(n9445), .A2(n10004), .B1(n9444), .B2(n10036), .ZN(n1376) );
  OAI221_X1 U1104 ( .B1(n8523), .B2(n9500), .C1(n8491), .C2(n9497), .A(n1224), 
        .ZN(n1219) );
  AOI22_X1 U1105 ( .A1(n9494), .A2(n10492), .B1(n9491), .B2(n10364), .ZN(n1224) );
  OAI221_X1 U1106 ( .B1(n8510), .B2(n9499), .C1(n8478), .C2(n9496), .A(n1465), 
        .ZN(n1453) );
  AOI22_X1 U1107 ( .A1(n9493), .A2(n10505), .B1(n9492), .B2(n10377), .ZN(n1465) );
  OAI221_X1 U1108 ( .B1(n8524), .B2(n9500), .C1(n8492), .C2(n9497), .A(n1206), 
        .ZN(n1201) );
  AOI22_X1 U1109 ( .A1(n9494), .A2(n10491), .B1(n9491), .B2(n10363), .ZN(n1206) );
  OAI221_X1 U1110 ( .B1(n8525), .B2(n9500), .C1(n8493), .C2(n9497), .A(n1188), 
        .ZN(n1183) );
  AOI22_X1 U1111 ( .A1(n9494), .A2(n10490), .B1(n9491), .B2(n10362), .ZN(n1188) );
  OAI221_X1 U1112 ( .B1(n8530), .B2(n9500), .C1(n8498), .C2(n9497), .A(n1098), 
        .ZN(n1093) );
  AOI22_X1 U1113 ( .A1(n9494), .A2(n10485), .B1(n9490), .B2(n10357), .ZN(n1098) );
  OAI221_X1 U1114 ( .B1(n8850), .B2(n9452), .C1(n8818), .C2(n9449), .A(n1106), 
        .ZN(n1101) );
  AOI22_X1 U1115 ( .A1(n9446), .A2(n9989), .B1(n9442), .B2(n10021), .ZN(n1106)
         );
  OAI221_X1 U1116 ( .B1(n8845), .B2(n9452), .C1(n8813), .C2(n9449), .A(n1196), 
        .ZN(n1191) );
  AOI22_X1 U1117 ( .A1(n9446), .A2(n9994), .B1(n9443), .B2(n10026), .ZN(n1196)
         );
  OAI221_X1 U1118 ( .B1(n8520), .B2(n9499), .C1(n8488), .C2(n9496), .A(n1278), 
        .ZN(n1273) );
  AOI22_X1 U1119 ( .A1(n9493), .A2(n10495), .B1(n9491), .B2(n10367), .ZN(n1278) );
  OAI221_X1 U1120 ( .B1(n8521), .B2(n9499), .C1(n8489), .C2(n9496), .A(n1260), 
        .ZN(n1255) );
  AOI22_X1 U1121 ( .A1(n9493), .A2(n10494), .B1(n9491), .B2(n10366), .ZN(n1260) );
  OAI221_X1 U1122 ( .B1(n8532), .B2(n9500), .C1(n8500), .C2(n9497), .A(n1062), 
        .ZN(n1057) );
  AOI22_X1 U1123 ( .A1(n9494), .A2(n10483), .B1(n9490), .B2(n10355), .ZN(n1062) );
  OAI221_X1 U1124 ( .B1(n8531), .B2(n9500), .C1(n8499), .C2(n9497), .A(n1080), 
        .ZN(n1075) );
  AOI22_X1 U1125 ( .A1(n9494), .A2(n10484), .B1(n9490), .B2(n10356), .ZN(n1080) );
  OAI221_X1 U1126 ( .B1(n8851), .B2(n9452), .C1(n8819), .C2(n9449), .A(n1088), 
        .ZN(n1083) );
  AOI22_X1 U1127 ( .A1(n9446), .A2(n9988), .B1(n9442), .B2(n10020), .ZN(n1088)
         );
  OAI221_X1 U1128 ( .B1(n8841), .B2(n9451), .C1(n8809), .C2(n9448), .A(n1268), 
        .ZN(n1263) );
  AOI22_X1 U1129 ( .A1(n9445), .A2(n9998), .B1(n9443), .B2(n10030), .ZN(n1268)
         );
  OAI221_X1 U1130 ( .B1(n8852), .B2(n9452), .C1(n8820), .C2(n9449), .A(n1070), 
        .ZN(n1065) );
  AOI22_X1 U1131 ( .A1(n9446), .A2(n9987), .B1(n9442), .B2(n10019), .ZN(n1070)
         );
  OAI221_X1 U1132 ( .B1(n8526), .B2(n9500), .C1(n8494), .C2(n9497), .A(n1170), 
        .ZN(n1165) );
  AOI22_X1 U1133 ( .A1(n9494), .A2(n10489), .B1(n9491), .B2(n10361), .ZN(n1170) );
  OAI221_X1 U1134 ( .B1(n8846), .B2(n9452), .C1(n8814), .C2(n9449), .A(n1178), 
        .ZN(n1173) );
  AOI22_X1 U1135 ( .A1(n9446), .A2(n9993), .B1(n9443), .B2(n10025), .ZN(n1178)
         );
  OAI221_X1 U1136 ( .B1(n8522), .B2(n9500), .C1(n8490), .C2(n9497), .A(n1242), 
        .ZN(n1237) );
  AOI22_X1 U1137 ( .A1(n9494), .A2(n10493), .B1(n9491), .B2(n10365), .ZN(n1242) );
  OAI221_X1 U1138 ( .B1(n8533), .B2(n9500), .C1(n8501), .C2(n9497), .A(n1044), 
        .ZN(n1039) );
  AOI22_X1 U1139 ( .A1(n9494), .A2(n10482), .B1(n9490), .B2(n10354), .ZN(n1044) );
  OAI221_X1 U1140 ( .B1(n8842), .B2(n9452), .C1(n8810), .C2(n9449), .A(n1250), 
        .ZN(n1245) );
  AOI22_X1 U1141 ( .A1(n9446), .A2(n9997), .B1(n9443), .B2(n10029), .ZN(n1250)
         );
  OAI221_X1 U1142 ( .B1(n8853), .B2(n9452), .C1(n8821), .C2(n9449), .A(n1052), 
        .ZN(n1047) );
  AOI22_X1 U1143 ( .A1(n9446), .A2(n9986), .B1(n9442), .B2(n10018), .ZN(n1052)
         );
  OAI221_X1 U1144 ( .B1(n8527), .B2(n9500), .C1(n8495), .C2(n9497), .A(n1152), 
        .ZN(n1147) );
  AOI22_X1 U1145 ( .A1(n9494), .A2(n10488), .B1(n9491), .B2(n10360), .ZN(n1152) );
  OAI221_X1 U1146 ( .B1(n8528), .B2(n9500), .C1(n8496), .C2(n9497), .A(n1134), 
        .ZN(n1129) );
  AOI22_X1 U1147 ( .A1(n9494), .A2(n10487), .B1(n9491), .B2(n10359), .ZN(n1134) );
  OAI221_X1 U1148 ( .B1(n8529), .B2(n9500), .C1(n8497), .C2(n9497), .A(n1116), 
        .ZN(n1111) );
  AOI22_X1 U1149 ( .A1(n9494), .A2(n10486), .B1(n9491), .B2(n10358), .ZN(n1116) );
  OAI221_X1 U1150 ( .B1(n8849), .B2(n9452), .C1(n8817), .C2(n9449), .A(n1124), 
        .ZN(n1119) );
  AOI22_X1 U1151 ( .A1(n9446), .A2(n9990), .B1(n9443), .B2(n10022), .ZN(n1124)
         );
  OAI221_X1 U1152 ( .B1(n8511), .B2(n9499), .C1(n8479), .C2(n9496), .A(n1440), 
        .ZN(n1435) );
  AOI22_X1 U1153 ( .A1(n9493), .A2(n10504), .B1(n9492), .B2(n10376), .ZN(n1440) );
  OAI221_X1 U1154 ( .B1(n8831), .B2(n9451), .C1(n8799), .C2(n9448), .A(n1448), 
        .ZN(n1443) );
  AOI22_X1 U1155 ( .A1(n9445), .A2(n10008), .B1(n9444), .B2(n10040), .ZN(n1448) );
  OAI221_X1 U1156 ( .B1(n8512), .B2(n9499), .C1(n8480), .C2(n9496), .A(n1422), 
        .ZN(n1417) );
  AOI22_X1 U1157 ( .A1(n9493), .A2(n10503), .B1(n9492), .B2(n10375), .ZN(n1422) );
  OAI221_X1 U1158 ( .B1(n8535), .B2(n9501), .C1(n8503), .C2(n9498), .A(n1008), 
        .ZN(n1003) );
  AOI22_X1 U1159 ( .A1(n9495), .A2(n10480), .B1(n9490), .B2(n10352), .ZN(n1008) );
  OAI221_X1 U1160 ( .B1(n8538), .B2(n9501), .C1(n8506), .C2(n9498), .A(n954), 
        .ZN(n949) );
  AOI22_X1 U1161 ( .A1(n9495), .A2(n10477), .B1(n9490), .B2(n10349), .ZN(n954)
         );
  OAI221_X1 U1162 ( .B1(n8855), .B2(n9453), .C1(n8823), .C2(n9450), .A(n1016), 
        .ZN(n1011) );
  AOI22_X1 U1163 ( .A1(n9447), .A2(n10576), .B1(n9442), .B2(n10016), .ZN(n1016) );
  OAI221_X1 U1164 ( .B1(n8516), .B2(n9499), .C1(n8484), .C2(n9496), .A(n1350), 
        .ZN(n1345) );
  AOI22_X1 U1165 ( .A1(n9493), .A2(n10499), .B1(n9492), .B2(n10371), .ZN(n1350) );
  OAI221_X1 U1166 ( .B1(n8832), .B2(n9451), .C1(n8800), .C2(n9448), .A(n1430), 
        .ZN(n1425) );
  AOI22_X1 U1167 ( .A1(n9445), .A2(n10007), .B1(n9444), .B2(n10039), .ZN(n1430) );
  OAI221_X1 U1168 ( .B1(n8534), .B2(n9501), .C1(n8502), .C2(n9498), .A(n1026), 
        .ZN(n1021) );
  AOI22_X1 U1169 ( .A1(n9495), .A2(n10481), .B1(n9490), .B2(n10353), .ZN(n1026) );
  OAI221_X1 U1170 ( .B1(n8539), .B2(n9501), .C1(n8507), .C2(n9498), .A(n936), 
        .ZN(n931) );
  AOI22_X1 U1171 ( .A1(n9495), .A2(n10476), .B1(n9490), .B2(n10348), .ZN(n936)
         );
  OAI221_X1 U1172 ( .B1(n8517), .B2(n9499), .C1(n8485), .C2(n9496), .A(n1332), 
        .ZN(n1327) );
  AOI22_X1 U1173 ( .A1(n9493), .A2(n10498), .B1(n9492), .B2(n10370), .ZN(n1332) );
  OAI221_X1 U1174 ( .B1(n8837), .B2(n9451), .C1(n8805), .C2(n9448), .A(n1340), 
        .ZN(n1335) );
  AOI22_X1 U1175 ( .A1(n9445), .A2(n10002), .B1(n9444), .B2(n10034), .ZN(n1340) );
  OAI221_X1 U1176 ( .B1(n8536), .B2(n9501), .C1(n8504), .C2(n9498), .A(n990), 
        .ZN(n985) );
  AOI22_X1 U1177 ( .A1(n9495), .A2(n10479), .B1(n9490), .B2(n10351), .ZN(n990)
         );
  OAI221_X1 U1178 ( .B1(n8856), .B2(n9453), .C1(n8824), .C2(n9450), .A(n998), 
        .ZN(n993) );
  AOI22_X1 U1179 ( .A1(n9447), .A2(n10575), .B1(n9442), .B2(n10015), .ZN(n998)
         );
  OAI221_X1 U1180 ( .B1(n8540), .B2(n9501), .C1(n8508), .C2(n9498), .A(n918), 
        .ZN(n913) );
  AOI22_X1 U1181 ( .A1(n9495), .A2(n10475), .B1(n9490), .B2(n10347), .ZN(n918)
         );
  OAI221_X1 U1182 ( .B1(n8518), .B2(n9499), .C1(n8486), .C2(n9496), .A(n1314), 
        .ZN(n1309) );
  AOI22_X1 U1183 ( .A1(n9493), .A2(n10497), .B1(n9491), .B2(n10369), .ZN(n1314) );
  OAI221_X1 U1184 ( .B1(n8838), .B2(n9451), .C1(n8806), .C2(n9448), .A(n1322), 
        .ZN(n1317) );
  AOI22_X1 U1185 ( .A1(n9445), .A2(n10001), .B1(n9443), .B2(n10033), .ZN(n1322) );
  OAI221_X1 U1186 ( .B1(n8860), .B2(n9453), .C1(n8828), .C2(n9450), .A(n926), 
        .ZN(n921) );
  AOI22_X1 U1187 ( .A1(n9447), .A2(n10571), .B1(n9442), .B2(n10011), .ZN(n926)
         );
  OAI221_X1 U1188 ( .B1(n8537), .B2(n9501), .C1(n8505), .C2(n9498), .A(n972), 
        .ZN(n967) );
  AOI22_X1 U1189 ( .A1(n9495), .A2(n10478), .B1(n9490), .B2(n10350), .ZN(n972)
         );
  OAI221_X1 U1190 ( .B1(n8519), .B2(n9499), .C1(n8487), .C2(n9496), .A(n1296), 
        .ZN(n1291) );
  AOI22_X1 U1191 ( .A1(n9493), .A2(n10496), .B1(n9491), .B2(n10368), .ZN(n1296) );
  OAI221_X1 U1192 ( .B1(n8857), .B2(n9453), .C1(n8825), .C2(n9450), .A(n980), 
        .ZN(n975) );
  AOI22_X1 U1193 ( .A1(n9447), .A2(n10574), .B1(n9442), .B2(n10014), .ZN(n980)
         );
  OAI221_X1 U1194 ( .B1(n8839), .B2(n9451), .C1(n8807), .C2(n9448), .A(n1304), 
        .ZN(n1299) );
  AOI22_X1 U1195 ( .A1(n9445), .A2(n10000), .B1(n9443), .B2(n10032), .ZN(n1304) );
  OAI221_X1 U1196 ( .B1(n8806), .B2(n9355), .C1(n8782), .C2(n9352), .A(n1942), 
        .ZN(n1937) );
  AOI22_X1 U1197 ( .A1(n9349), .A2(n10033), .B1(n9347), .B2(n10065), .ZN(n1942) );
  OAI221_X1 U1198 ( .B1(n8807), .B2(n9355), .C1(n8783), .C2(n9352), .A(n1924), 
        .ZN(n1919) );
  AOI22_X1 U1199 ( .A1(n9349), .A2(n10032), .B1(n9347), .B2(n10064), .ZN(n1924) );
  OAI221_X1 U1200 ( .B1(n8808), .B2(n9355), .C1(n8784), .C2(n9352), .A(n1906), 
        .ZN(n1901) );
  AOI22_X1 U1201 ( .A1(n9349), .A2(n10031), .B1(n9347), .B2(n10063), .ZN(n1906) );
  OAI221_X1 U1202 ( .B1(n8809), .B2(n9355), .C1(n8785), .C2(n9352), .A(n1888), 
        .ZN(n1883) );
  AOI22_X1 U1203 ( .A1(n9349), .A2(n10030), .B1(n9347), .B2(n10062), .ZN(n1888) );
  OAI221_X1 U1204 ( .B1(n8810), .B2(n9356), .C1(n8786), .C2(n9353), .A(n1870), 
        .ZN(n1865) );
  AOI22_X1 U1205 ( .A1(n9350), .A2(n10029), .B1(n9347), .B2(n10061), .ZN(n1870) );
  OAI221_X1 U1206 ( .B1(n8811), .B2(n9356), .C1(n8787), .C2(n9353), .A(n1852), 
        .ZN(n1847) );
  AOI22_X1 U1207 ( .A1(n9350), .A2(n10028), .B1(n9347), .B2(n10060), .ZN(n1852) );
  OAI221_X1 U1208 ( .B1(n8812), .B2(n9356), .C1(n8788), .C2(n9353), .A(n1834), 
        .ZN(n1829) );
  AOI22_X1 U1209 ( .A1(n9350), .A2(n10027), .B1(n9347), .B2(n10059), .ZN(n1834) );
  OAI221_X1 U1210 ( .B1(n8813), .B2(n9356), .C1(n8789), .C2(n9353), .A(n1816), 
        .ZN(n1811) );
  AOI22_X1 U1211 ( .A1(n9350), .A2(n10026), .B1(n9347), .B2(n10058), .ZN(n1816) );
  OAI221_X1 U1212 ( .B1(n8814), .B2(n9356), .C1(n8790), .C2(n9353), .A(n1798), 
        .ZN(n1793) );
  AOI22_X1 U1213 ( .A1(n9350), .A2(n10025), .B1(n9347), .B2(n10057), .ZN(n1798) );
  OAI221_X1 U1214 ( .B1(n8815), .B2(n9356), .C1(n8791), .C2(n9353), .A(n1780), 
        .ZN(n1775) );
  AOI22_X1 U1215 ( .A1(n9350), .A2(n10024), .B1(n9347), .B2(n10056), .ZN(n1780) );
  OAI221_X1 U1216 ( .B1(n8816), .B2(n9356), .C1(n8792), .C2(n9353), .A(n1762), 
        .ZN(n1757) );
  AOI22_X1 U1217 ( .A1(n9350), .A2(n10023), .B1(n9347), .B2(n10055), .ZN(n1762) );
  OAI221_X1 U1218 ( .B1(n8817), .B2(n9356), .C1(n8793), .C2(n9353), .A(n1744), 
        .ZN(n1739) );
  AOI22_X1 U1219 ( .A1(n9350), .A2(n10022), .B1(n9347), .B2(n10054), .ZN(n1744) );
  OAI221_X1 U1220 ( .B1(n8818), .B2(n9356), .C1(n8794), .C2(n9353), .A(n1726), 
        .ZN(n1721) );
  AOI22_X1 U1221 ( .A1(n9350), .A2(n10021), .B1(n9346), .B2(n10053), .ZN(n1726) );
  OAI221_X1 U1222 ( .B1(n8819), .B2(n9356), .C1(n8795), .C2(n9353), .A(n1708), 
        .ZN(n1703) );
  AOI22_X1 U1223 ( .A1(n9350), .A2(n10020), .B1(n9346), .B2(n10052), .ZN(n1708) );
  OAI221_X1 U1224 ( .B1(n8820), .B2(n9356), .C1(n8796), .C2(n9353), .A(n1690), 
        .ZN(n1685) );
  AOI22_X1 U1225 ( .A1(n9350), .A2(n10019), .B1(n9346), .B2(n10051), .ZN(n1690) );
  OAI221_X1 U1226 ( .B1(n8821), .B2(n9356), .C1(n8797), .C2(n9353), .A(n1672), 
        .ZN(n1667) );
  AOI22_X1 U1227 ( .A1(n9350), .A2(n10018), .B1(n9346), .B2(n10050), .ZN(n1672) );
  OAI221_X1 U1228 ( .B1(n8822), .B2(n9357), .C1(n8311), .C2(n9354), .A(n1654), 
        .ZN(n1649) );
  AOI22_X1 U1229 ( .A1(n9351), .A2(n10017), .B1(n9346), .B2(n10049), .ZN(n1654) );
  OAI221_X1 U1230 ( .B1(n8823), .B2(n9357), .C1(n8312), .C2(n9354), .A(n1636), 
        .ZN(n1631) );
  AOI22_X1 U1231 ( .A1(n9351), .A2(n10016), .B1(n9346), .B2(n10048), .ZN(n1636) );
  OAI221_X1 U1232 ( .B1(n8824), .B2(n9357), .C1(n8313), .C2(n9354), .A(n1618), 
        .ZN(n1613) );
  AOI22_X1 U1233 ( .A1(n9351), .A2(n10015), .B1(n9346), .B2(n10047), .ZN(n1618) );
  OAI221_X1 U1234 ( .B1(n8825), .B2(n9357), .C1(n8314), .C2(n9354), .A(n1600), 
        .ZN(n1595) );
  AOI22_X1 U1235 ( .A1(n9351), .A2(n10014), .B1(n9346), .B2(n10046), .ZN(n1600) );
  OAI221_X1 U1236 ( .B1(n8826), .B2(n9357), .C1(n8315), .C2(n9354), .A(n1582), 
        .ZN(n1577) );
  AOI22_X1 U1237 ( .A1(n9351), .A2(n10013), .B1(n9346), .B2(n10045), .ZN(n1582) );
  OAI221_X1 U1238 ( .B1(n8827), .B2(n9357), .C1(n8316), .C2(n9354), .A(n1564), 
        .ZN(n1559) );
  AOI22_X1 U1239 ( .A1(n9351), .A2(n10012), .B1(n9346), .B2(n10044), .ZN(n1564) );
  OAI221_X1 U1240 ( .B1(n8828), .B2(n9357), .C1(n8317), .C2(n9354), .A(n1546), 
        .ZN(n1541) );
  AOI22_X1 U1241 ( .A1(n9351), .A2(n10011), .B1(n9346), .B2(n10043), .ZN(n1546) );
  OAI221_X1 U1242 ( .B1(n8829), .B2(n9357), .C1(n8318), .C2(n9354), .A(n1522), 
        .ZN(n1507) );
  AOI22_X1 U1243 ( .A1(n9351), .A2(n10010), .B1(n9346), .B2(n10042), .ZN(n1522) );
  OAI221_X1 U1244 ( .B1(n8922), .B2(n9439), .C1(n8890), .C2(n9436), .A(n1395), 
        .ZN(n1388) );
  AOI22_X1 U1245 ( .A1(n9433), .A2(n10341), .B1(n9432), .B2(n9949), .ZN(n1395)
         );
  OAI221_X1 U1246 ( .B1(n8923), .B2(n9439), .C1(n8891), .C2(n9436), .A(n1377), 
        .ZN(n1370) );
  AOI22_X1 U1247 ( .A1(n9433), .A2(n10340), .B1(n9432), .B2(n9948), .ZN(n1377)
         );
  OAI221_X1 U1248 ( .B1(n2247), .B2(n9488), .C1(n8388), .C2(n9485), .A(n1225), 
        .ZN(n1218) );
  AOI22_X1 U1249 ( .A1(n9482), .A2(n10212), .B1(n9479), .B2(n10644), .ZN(n1225) );
  OAI221_X1 U1250 ( .B1(n2239), .B2(n9488), .C1(n8389), .C2(n9485), .A(n1207), 
        .ZN(n1200) );
  AOI22_X1 U1251 ( .A1(n9482), .A2(n10211), .B1(n9479), .B2(n10643), .ZN(n1207) );
  OAI221_X1 U1252 ( .B1(n2231), .B2(n9488), .C1(n8390), .C2(n9485), .A(n1189), 
        .ZN(n1182) );
  AOI22_X1 U1253 ( .A1(n9482), .A2(n10210), .B1(n9479), .B2(n10642), .ZN(n1189) );
  OAI221_X1 U1254 ( .B1(n2191), .B2(n9488), .C1(n8395), .C2(n9485), .A(n1099), 
        .ZN(n1092) );
  AOI22_X1 U1255 ( .A1(n9482), .A2(n10205), .B1(n9478), .B2(n10637), .ZN(n1099) );
  OAI221_X1 U1256 ( .B1(n2271), .B2(n9487), .C1(n8385), .C2(n9484), .A(n1279), 
        .ZN(n1272) );
  AOI22_X1 U1257 ( .A1(n9481), .A2(n10215), .B1(n9479), .B2(n10647), .ZN(n1279) );
  OAI221_X1 U1258 ( .B1(n2263), .B2(n9487), .C1(n8386), .C2(n9484), .A(n1261), 
        .ZN(n1254) );
  AOI22_X1 U1259 ( .A1(n9481), .A2(n10214), .B1(n9479), .B2(n10646), .ZN(n1261) );
  OAI221_X1 U1260 ( .B1(n2175), .B2(n9488), .C1(n8397), .C2(n9485), .A(n1063), 
        .ZN(n1056) );
  AOI22_X1 U1261 ( .A1(n9482), .A2(n10203), .B1(n9478), .B2(n10635), .ZN(n1063) );
  OAI221_X1 U1262 ( .B1(n2183), .B2(n9488), .C1(n8396), .C2(n9485), .A(n1081), 
        .ZN(n1074) );
  AOI22_X1 U1263 ( .A1(n9482), .A2(n10204), .B1(n9478), .B2(n10636), .ZN(n1081) );
  OAI221_X1 U1264 ( .B1(n8938), .B2(n9440), .C1(n8906), .C2(n9437), .A(n1107), 
        .ZN(n1100) );
  AOI22_X1 U1265 ( .A1(n9434), .A2(n10325), .B1(n9430), .B2(n9933), .ZN(n1107)
         );
  OAI221_X1 U1266 ( .B1(n8933), .B2(n9440), .C1(n8901), .C2(n9437), .A(n1197), 
        .ZN(n1190) );
  AOI22_X1 U1267 ( .A1(n9434), .A2(n10330), .B1(n9431), .B2(n9938), .ZN(n1197)
         );
  OAI221_X1 U1268 ( .B1(n8939), .B2(n9440), .C1(n8907), .C2(n9437), .A(n1089), 
        .ZN(n1082) );
  AOI22_X1 U1269 ( .A1(n9434), .A2(n10324), .B1(n9430), .B2(n9932), .ZN(n1089)
         );
  OAI221_X1 U1270 ( .B1(n8929), .B2(n9439), .C1(n8897), .C2(n9436), .A(n1269), 
        .ZN(n1262) );
  AOI22_X1 U1271 ( .A1(n9433), .A2(n10334), .B1(n9431), .B2(n9942), .ZN(n1269)
         );
  OAI221_X1 U1272 ( .B1(n8940), .B2(n9440), .C1(n8908), .C2(n9437), .A(n1071), 
        .ZN(n1064) );
  AOI22_X1 U1273 ( .A1(n9434), .A2(n10323), .B1(n9430), .B2(n9931), .ZN(n1071)
         );
  OAI221_X1 U1274 ( .B1(n2223), .B2(n9488), .C1(n8391), .C2(n9485), .A(n1171), 
        .ZN(n1164) );
  AOI22_X1 U1275 ( .A1(n9482), .A2(n10209), .B1(n9479), .B2(n10641), .ZN(n1171) );
  OAI221_X1 U1276 ( .B1(n2255), .B2(n9488), .C1(n8387), .C2(n9485), .A(n1243), 
        .ZN(n1236) );
  AOI22_X1 U1277 ( .A1(n9482), .A2(n10213), .B1(n9479), .B2(n10645), .ZN(n1243) );
  OAI221_X1 U1278 ( .B1(n2167), .B2(n9488), .C1(n8398), .C2(n9485), .A(n1045), 
        .ZN(n1038) );
  AOI22_X1 U1279 ( .A1(n9482), .A2(n10202), .B1(n9478), .B2(n10634), .ZN(n1045) );
  OAI221_X1 U1280 ( .B1(n8934), .B2(n9440), .C1(n8902), .C2(n9437), .A(n1179), 
        .ZN(n1172) );
  AOI22_X1 U1281 ( .A1(n9434), .A2(n10329), .B1(n9431), .B2(n9937), .ZN(n1179)
         );
  OAI221_X1 U1282 ( .B1(n8930), .B2(n9440), .C1(n8898), .C2(n9437), .A(n1251), 
        .ZN(n1244) );
  AOI22_X1 U1283 ( .A1(n9434), .A2(n10333), .B1(n9431), .B2(n9941), .ZN(n1251)
         );
  OAI221_X1 U1284 ( .B1(n8941), .B2(n9440), .C1(n8909), .C2(n9437), .A(n1053), 
        .ZN(n1046) );
  AOI22_X1 U1285 ( .A1(n9434), .A2(n10322), .B1(n9430), .B2(n9930), .ZN(n1053)
         );
  OAI221_X1 U1286 ( .B1(n2215), .B2(n9488), .C1(n8392), .C2(n9485), .A(n1153), 
        .ZN(n1146) );
  AOI22_X1 U1287 ( .A1(n9482), .A2(n10208), .B1(n9479), .B2(n10640), .ZN(n1153) );
  OAI221_X1 U1288 ( .B1(n2207), .B2(n9488), .C1(n8393), .C2(n9485), .A(n1135), 
        .ZN(n1128) );
  AOI22_X1 U1289 ( .A1(n9482), .A2(n10207), .B1(n9479), .B2(n10639), .ZN(n1135) );
  OAI221_X1 U1290 ( .B1(n2199), .B2(n9488), .C1(n8394), .C2(n9485), .A(n1117), 
        .ZN(n1110) );
  AOI22_X1 U1291 ( .A1(n9482), .A2(n10206), .B1(n9479), .B2(n10638), .ZN(n1117) );
  OAI221_X1 U1292 ( .B1(n8937), .B2(n9440), .C1(n8905), .C2(n9437), .A(n1125), 
        .ZN(n1118) );
  AOI22_X1 U1293 ( .A1(n9434), .A2(n10326), .B1(n9431), .B2(n9934), .ZN(n1125)
         );
  OAI221_X1 U1294 ( .B1(n8919), .B2(n9439), .C1(n8887), .C2(n9436), .A(n1449), 
        .ZN(n1442) );
  AOI22_X1 U1295 ( .A1(n9433), .A2(n10344), .B1(n9432), .B2(n9952), .ZN(n1449)
         );
  OAI221_X1 U1296 ( .B1(n8920), .B2(n9439), .C1(n8888), .C2(n9436), .A(n1431), 
        .ZN(n1424) );
  AOI22_X1 U1297 ( .A1(n9433), .A2(n10343), .B1(n9432), .B2(n9951), .ZN(n1431)
         );
  OAI221_X1 U1298 ( .B1(n8943), .B2(n9441), .C1(n8911), .C2(n9438), .A(n1017), 
        .ZN(n1010) );
  AOI22_X1 U1299 ( .A1(n9435), .A2(n10568), .B1(n9430), .B2(n9928), .ZN(n1017)
         );
  OAI221_X1 U1300 ( .B1(n8925), .B2(n9439), .C1(n8893), .C2(n9436), .A(n1341), 
        .ZN(n1334) );
  AOI22_X1 U1301 ( .A1(n9433), .A2(n10338), .B1(n9432), .B2(n9946), .ZN(n1341)
         );
  OAI221_X1 U1302 ( .B1(n2287), .B2(n9487), .C1(n8383), .C2(n9484), .A(n1315), 
        .ZN(n1308) );
  AOI22_X1 U1303 ( .A1(n9481), .A2(n10217), .B1(n9479), .B2(n10649), .ZN(n1315) );
  OAI221_X1 U1304 ( .B1(n8944), .B2(n9441), .C1(n8912), .C2(n9438), .A(n999), 
        .ZN(n992) );
  AOI22_X1 U1305 ( .A1(n9435), .A2(n10567), .B1(n9430), .B2(n9927), .ZN(n999)
         );
  OAI221_X1 U1306 ( .B1(n2279), .B2(n9487), .C1(n8384), .C2(n9484), .A(n1297), 
        .ZN(n1290) );
  AOI22_X1 U1307 ( .A1(n9481), .A2(n10216), .B1(n9479), .B2(n10648), .ZN(n1297) );
  OAI221_X1 U1308 ( .B1(n8926), .B2(n9439), .C1(n8894), .C2(n9436), .A(n1323), 
        .ZN(n1316) );
  AOI22_X1 U1309 ( .A1(n9433), .A2(n10337), .B1(n9431), .B2(n9945), .ZN(n1323)
         );
  OAI221_X1 U1310 ( .B1(n8948), .B2(n9441), .C1(n8916), .C2(n9438), .A(n927), 
        .ZN(n920) );
  AOI22_X1 U1311 ( .A1(n9435), .A2(n10563), .B1(n9430), .B2(n9923), .ZN(n927)
         );
  OAI221_X1 U1312 ( .B1(n8945), .B2(n9441), .C1(n8913), .C2(n9438), .A(n981), 
        .ZN(n974) );
  AOI22_X1 U1313 ( .A1(n9435), .A2(n10566), .B1(n9430), .B2(n9926), .ZN(n981)
         );
  OAI221_X1 U1314 ( .B1(n8927), .B2(n9439), .C1(n8895), .C2(n9436), .A(n1305), 
        .ZN(n1298) );
  AOI22_X1 U1315 ( .A1(n9433), .A2(n10336), .B1(n9431), .B2(n9944), .ZN(n1305)
         );
  OAI221_X1 U1316 ( .B1(n8894), .B2(n9343), .C1(n8870), .C2(n9340), .A(n1943), 
        .ZN(n1936) );
  AOI22_X1 U1317 ( .A1(n9337), .A2(n9945), .B1(n9335), .B2(n9977), .ZN(n1943)
         );
  OAI221_X1 U1318 ( .B1(n8895), .B2(n9343), .C1(n8871), .C2(n9340), .A(n1925), 
        .ZN(n1918) );
  AOI22_X1 U1319 ( .A1(n9337), .A2(n9944), .B1(n9335), .B2(n9976), .ZN(n1925)
         );
  OAI221_X1 U1320 ( .B1(n8896), .B2(n9343), .C1(n8872), .C2(n9340), .A(n1907), 
        .ZN(n1900) );
  AOI22_X1 U1321 ( .A1(n9337), .A2(n9943), .B1(n9335), .B2(n9975), .ZN(n1907)
         );
  OAI221_X1 U1322 ( .B1(n8897), .B2(n9343), .C1(n8873), .C2(n9340), .A(n1889), 
        .ZN(n1882) );
  AOI22_X1 U1323 ( .A1(n9337), .A2(n9942), .B1(n9335), .B2(n9974), .ZN(n1889)
         );
  OAI221_X1 U1324 ( .B1(n8898), .B2(n9344), .C1(n8874), .C2(n9341), .A(n1871), 
        .ZN(n1864) );
  AOI22_X1 U1325 ( .A1(n9338), .A2(n9941), .B1(n9335), .B2(n9973), .ZN(n1871)
         );
  OAI221_X1 U1326 ( .B1(n8899), .B2(n9344), .C1(n8875), .C2(n9341), .A(n1853), 
        .ZN(n1846) );
  AOI22_X1 U1327 ( .A1(n9338), .A2(n9940), .B1(n9335), .B2(n9972), .ZN(n1853)
         );
  OAI221_X1 U1328 ( .B1(n8900), .B2(n9344), .C1(n8876), .C2(n9341), .A(n1835), 
        .ZN(n1828) );
  AOI22_X1 U1329 ( .A1(n9338), .A2(n9939), .B1(n9335), .B2(n9971), .ZN(n1835)
         );
  OAI221_X1 U1330 ( .B1(n8901), .B2(n9344), .C1(n8877), .C2(n9341), .A(n1817), 
        .ZN(n1810) );
  AOI22_X1 U1331 ( .A1(n9338), .A2(n9938), .B1(n9335), .B2(n9970), .ZN(n1817)
         );
  OAI221_X1 U1332 ( .B1(n8902), .B2(n9344), .C1(n8878), .C2(n9341), .A(n1799), 
        .ZN(n1792) );
  AOI22_X1 U1333 ( .A1(n9338), .A2(n9937), .B1(n9335), .B2(n9969), .ZN(n1799)
         );
  OAI221_X1 U1334 ( .B1(n8903), .B2(n9344), .C1(n8879), .C2(n9341), .A(n1781), 
        .ZN(n1774) );
  AOI22_X1 U1335 ( .A1(n9338), .A2(n9936), .B1(n9335), .B2(n9968), .ZN(n1781)
         );
  OAI221_X1 U1336 ( .B1(n8904), .B2(n9344), .C1(n8880), .C2(n9341), .A(n1763), 
        .ZN(n1756) );
  AOI22_X1 U1337 ( .A1(n9338), .A2(n9935), .B1(n9335), .B2(n9967), .ZN(n1763)
         );
  OAI221_X1 U1338 ( .B1(n8905), .B2(n9344), .C1(n8881), .C2(n9341), .A(n1745), 
        .ZN(n1738) );
  AOI22_X1 U1339 ( .A1(n9338), .A2(n9934), .B1(n9335), .B2(n9966), .ZN(n1745)
         );
  OAI221_X1 U1340 ( .B1(n8906), .B2(n9344), .C1(n8882), .C2(n9341), .A(n1727), 
        .ZN(n1720) );
  AOI22_X1 U1341 ( .A1(n9338), .A2(n9933), .B1(n9334), .B2(n9965), .ZN(n1727)
         );
  OAI221_X1 U1342 ( .B1(n8907), .B2(n9344), .C1(n8883), .C2(n9341), .A(n1709), 
        .ZN(n1702) );
  AOI22_X1 U1343 ( .A1(n9338), .A2(n9932), .B1(n9334), .B2(n9964), .ZN(n1709)
         );
  OAI221_X1 U1344 ( .B1(n8908), .B2(n9344), .C1(n8884), .C2(n9341), .A(n1691), 
        .ZN(n1684) );
  AOI22_X1 U1345 ( .A1(n9338), .A2(n9931), .B1(n9334), .B2(n9963), .ZN(n1691)
         );
  OAI221_X1 U1346 ( .B1(n8909), .B2(n9344), .C1(n8885), .C2(n9341), .A(n1673), 
        .ZN(n1666) );
  AOI22_X1 U1347 ( .A1(n9338), .A2(n9930), .B1(n9334), .B2(n9962), .ZN(n1673)
         );
  OAI221_X1 U1348 ( .B1(n8910), .B2(n9345), .C1(n8303), .C2(n9342), .A(n1655), 
        .ZN(n1648) );
  AOI22_X1 U1349 ( .A1(n9339), .A2(n9929), .B1(n9334), .B2(n9961), .ZN(n1655)
         );
  OAI221_X1 U1350 ( .B1(n8911), .B2(n9345), .C1(n8304), .C2(n9342), .A(n1637), 
        .ZN(n1630) );
  AOI22_X1 U1351 ( .A1(n9339), .A2(n9928), .B1(n9334), .B2(n9960), .ZN(n1637)
         );
  OAI221_X1 U1352 ( .B1(n8912), .B2(n9345), .C1(n8305), .C2(n9342), .A(n1619), 
        .ZN(n1612) );
  AOI22_X1 U1353 ( .A1(n9339), .A2(n9927), .B1(n9334), .B2(n9959), .ZN(n1619)
         );
  OAI221_X1 U1354 ( .B1(n8913), .B2(n9345), .C1(n8306), .C2(n9342), .A(n1601), 
        .ZN(n1594) );
  AOI22_X1 U1355 ( .A1(n9339), .A2(n9926), .B1(n9334), .B2(n9958), .ZN(n1601)
         );
  OAI221_X1 U1356 ( .B1(n8914), .B2(n9345), .C1(n8307), .C2(n9342), .A(n1583), 
        .ZN(n1576) );
  AOI22_X1 U1357 ( .A1(n9339), .A2(n9925), .B1(n9334), .B2(n9957), .ZN(n1583)
         );
  OAI221_X1 U1358 ( .B1(n8915), .B2(n9345), .C1(n8308), .C2(n9342), .A(n1565), 
        .ZN(n1558) );
  AOI22_X1 U1359 ( .A1(n9339), .A2(n9924), .B1(n9334), .B2(n9956), .ZN(n1565)
         );
  OAI221_X1 U1360 ( .B1(n8916), .B2(n9345), .C1(n8309), .C2(n9342), .A(n1547), 
        .ZN(n1540) );
  AOI22_X1 U1361 ( .A1(n9339), .A2(n9923), .B1(n9334), .B2(n9955), .ZN(n1547)
         );
  OAI221_X1 U1362 ( .B1(n8917), .B2(n9345), .C1(n8310), .C2(n9342), .A(n1527), 
        .ZN(n1506) );
  AOI22_X1 U1363 ( .A1(n9339), .A2(n9922), .B1(n9334), .B2(n9954), .ZN(n1527)
         );
  AOI22_X1 U1364 ( .A1(n9458), .A2(n10124), .B1(n9455), .B2(n10156), .ZN(n1231) );
  AOI22_X1 U1365 ( .A1(n9457), .A2(n10137), .B1(n9456), .B2(n10169), .ZN(n1476) );
  AOI22_X1 U1366 ( .A1(n9458), .A2(n10120), .B1(n9455), .B2(n10152), .ZN(n1159) );
  AOI22_X1 U1367 ( .A1(n9457), .A2(n10131), .B1(n9456), .B2(n10163), .ZN(n1357) );
  AOI22_X1 U1368 ( .A1(n9470), .A2(n10180), .B1(n9467), .B2(n10244), .ZN(n1230) );
  AOI22_X1 U1369 ( .A1(n9469), .A2(n10193), .B1(n9468), .B2(n10257), .ZN(n1475) );
  AOI22_X1 U1370 ( .A1(n9470), .A2(n10176), .B1(n9467), .B2(n10240), .ZN(n1158) );
  AOI22_X1 U1371 ( .A1(n9469), .A2(n10187), .B1(n9468), .B2(n10251), .ZN(n1356) );
  NOR4_X1 U1372 ( .A1(n1452), .A2(n1453), .A3(n1454), .A4(n1455), .ZN(n1451)
         );
  OAI221_X1 U1373 ( .B1(n8918), .B2(n9439), .C1(n8886), .C2(n9436), .A(n1479), 
        .ZN(n1471) );
  NOR4_X1 U1374 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1217)
         );
  OAI221_X1 U1375 ( .B1(n8931), .B2(n9440), .C1(n8899), .C2(n9437), .A(n1233), 
        .ZN(n1226) );
  NOR4_X1 U1376 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1145)
         );
  OAI221_X1 U1377 ( .B1(n8935), .B2(n9440), .C1(n8903), .C2(n9437), .A(n1161), 
        .ZN(n1154) );
  NOR4_X1 U1378 ( .A1(n1308), .A2(n1309), .A3(n1310), .A4(n1311), .ZN(n1307)
         );
  NOR4_X1 U1379 ( .A1(n1316), .A2(n1317), .A3(n1318), .A4(n1319), .ZN(n1306)
         );
  OAI221_X1 U1380 ( .B1(n8247), .B2(n9511), .C1(n8228), .C2(n9508), .A(n1313), 
        .ZN(n1310) );
  OAI221_X1 U1381 ( .B1(n8921), .B2(n9439), .C1(n8889), .C2(n9436), .A(n1413), 
        .ZN(n1406) );
  AOI22_X1 U1382 ( .A1(n9433), .A2(n10342), .B1(n9432), .B2(n9950), .ZN(n1413)
         );
  OAI221_X1 U1383 ( .B1(n8949), .B2(n9441), .C1(n8917), .C2(n9438), .A(n907), 
        .ZN(n886) );
  AOI22_X1 U1384 ( .A1(n9435), .A2(n10562), .B1(n9430), .B2(n9922), .ZN(n907)
         );
  OAI221_X1 U1385 ( .B1(n8932), .B2(n9440), .C1(n8900), .C2(n9437), .A(n1215), 
        .ZN(n1208) );
  AOI22_X1 U1386 ( .A1(n9434), .A2(n10331), .B1(n9431), .B2(n9939), .ZN(n1215)
         );
  OAI221_X1 U1387 ( .B1(n8928), .B2(n9439), .C1(n8896), .C2(n9436), .A(n1287), 
        .ZN(n1280) );
  AOI22_X1 U1388 ( .A1(n9433), .A2(n10335), .B1(n9431), .B2(n9943), .ZN(n1287)
         );
  OAI221_X1 U1389 ( .B1(n8936), .B2(n9440), .C1(n8904), .C2(n9437), .A(n1143), 
        .ZN(n1136) );
  AOI22_X1 U1390 ( .A1(n9434), .A2(n10327), .B1(n9431), .B2(n9935), .ZN(n1143)
         );
  OAI221_X1 U1391 ( .B1(n8946), .B2(n9441), .C1(n8914), .C2(n9438), .A(n963), 
        .ZN(n956) );
  AOI22_X1 U1392 ( .A1(n9435), .A2(n10565), .B1(n9430), .B2(n9925), .ZN(n963)
         );
  OAI221_X1 U1393 ( .B1(n8942), .B2(n9441), .C1(n8910), .C2(n9438), .A(n1035), 
        .ZN(n1028) );
  AOI22_X1 U1394 ( .A1(n9435), .A2(n10569), .B1(n9430), .B2(n9929), .ZN(n1035)
         );
  OAI221_X1 U1395 ( .B1(n8947), .B2(n9441), .C1(n8915), .C2(n9438), .A(n945), 
        .ZN(n938) );
  AOI22_X1 U1396 ( .A1(n9435), .A2(n10564), .B1(n9430), .B2(n9924), .ZN(n945)
         );
  AND3_X1 U1397 ( .A1(ADD_RD2[4]), .A2(n10662), .A3(RD2), .ZN(n2088) );
  OAI221_X1 U1398 ( .B1(n8833), .B2(n9451), .C1(n8801), .C2(n9448), .A(n1412), 
        .ZN(n1407) );
  AOI22_X1 U1399 ( .A1(n9445), .A2(n10006), .B1(n9444), .B2(n10038), .ZN(n1412) );
  OAI221_X1 U1400 ( .B1(n8861), .B2(n9453), .C1(n8829), .C2(n9450), .A(n902), 
        .ZN(n887) );
  AOI22_X1 U1401 ( .A1(n9447), .A2(n10570), .B1(n9442), .B2(n10010), .ZN(n902)
         );
  OAI221_X1 U1402 ( .B1(n8843), .B2(n9452), .C1(n8811), .C2(n9449), .A(n1232), 
        .ZN(n1227) );
  AOI22_X1 U1403 ( .A1(n9446), .A2(n9996), .B1(n9443), .B2(n10028), .ZN(n1232)
         );
  OAI221_X1 U1404 ( .B1(n8830), .B2(n9451), .C1(n8798), .C2(n9448), .A(n1478), 
        .ZN(n1472) );
  AOI22_X1 U1405 ( .A1(n9445), .A2(n10009), .B1(n9444), .B2(n10041), .ZN(n1478) );
  OAI221_X1 U1406 ( .B1(n8844), .B2(n9452), .C1(n8812), .C2(n9449), .A(n1214), 
        .ZN(n1209) );
  AOI22_X1 U1407 ( .A1(n9446), .A2(n9995), .B1(n9443), .B2(n10027), .ZN(n1214)
         );
  OAI221_X1 U1408 ( .B1(n8840), .B2(n9451), .C1(n8808), .C2(n9448), .A(n1286), 
        .ZN(n1281) );
  AOI22_X1 U1409 ( .A1(n9445), .A2(n9999), .B1(n9443), .B2(n10031), .ZN(n1286)
         );
  OAI221_X1 U1410 ( .B1(n8847), .B2(n9452), .C1(n8815), .C2(n9449), .A(n1160), 
        .ZN(n1155) );
  AOI22_X1 U1411 ( .A1(n9446), .A2(n9992), .B1(n9443), .B2(n10024), .ZN(n1160)
         );
  OAI221_X1 U1412 ( .B1(n8848), .B2(n9452), .C1(n8816), .C2(n9449), .A(n1142), 
        .ZN(n1137) );
  AOI22_X1 U1413 ( .A1(n9446), .A2(n9991), .B1(n9443), .B2(n10023), .ZN(n1142)
         );
  OAI221_X1 U1414 ( .B1(n8858), .B2(n9453), .C1(n8826), .C2(n9450), .A(n962), 
        .ZN(n957) );
  AOI22_X1 U1415 ( .A1(n9447), .A2(n10573), .B1(n9442), .B2(n10013), .ZN(n962)
         );
  OAI221_X1 U1416 ( .B1(n8836), .B2(n9451), .C1(n8804), .C2(n9448), .A(n1358), 
        .ZN(n1353) );
  AOI22_X1 U1417 ( .A1(n9445), .A2(n10003), .B1(n9444), .B2(n10035), .ZN(n1358) );
  OAI221_X1 U1418 ( .B1(n8854), .B2(n9453), .C1(n8822), .C2(n9450), .A(n1034), 
        .ZN(n1029) );
  AOI22_X1 U1419 ( .A1(n9447), .A2(n10577), .B1(n9442), .B2(n10017), .ZN(n1034) );
  OAI221_X1 U1420 ( .B1(n8859), .B2(n9453), .C1(n8827), .C2(n9450), .A(n944), 
        .ZN(n939) );
  AOI22_X1 U1421 ( .A1(n9447), .A2(n10572), .B1(n9442), .B2(n10012), .ZN(n944)
         );
  OAI221_X1 U1422 ( .B1(n8777), .B2(n9463), .C1(n8239), .C2(n9460), .A(n1411), 
        .ZN(n1408) );
  AOI22_X1 U1423 ( .A1(n9457), .A2(n10134), .B1(n9456), .B2(n10166), .ZN(n1411) );
  OAI221_X1 U1424 ( .B1(n8318), .B2(n9465), .C1(n8183), .C2(n9462), .A(n897), 
        .ZN(n888) );
  AOI22_X1 U1425 ( .A1(n9459), .A2(n10106), .B1(n9454), .B2(n10138), .ZN(n897)
         );
  OAI221_X1 U1426 ( .B1(n8788), .B2(n9464), .C1(n8217), .C2(n9461), .A(n1213), 
        .ZN(n1210) );
  AOI22_X1 U1427 ( .A1(n9458), .A2(n10123), .B1(n9455), .B2(n10155), .ZN(n1213) );
  OAI221_X1 U1428 ( .B1(n8784), .B2(n9463), .C1(n8225), .C2(n9460), .A(n1285), 
        .ZN(n1282) );
  AOI22_X1 U1429 ( .A1(n9457), .A2(n10127), .B1(n9455), .B2(n10159), .ZN(n1285) );
  OAI221_X1 U1430 ( .B1(n8792), .B2(n9464), .C1(n8209), .C2(n9461), .A(n1141), 
        .ZN(n1138) );
  AOI22_X1 U1431 ( .A1(n9458), .A2(n10119), .B1(n9455), .B2(n10151), .ZN(n1141) );
  OAI221_X1 U1432 ( .B1(n8315), .B2(n9465), .C1(n8189), .C2(n9462), .A(n961), 
        .ZN(n958) );
  AOI22_X1 U1433 ( .A1(n9459), .A2(n10109), .B1(n9454), .B2(n10141), .ZN(n961)
         );
  OAI221_X1 U1434 ( .B1(n8311), .B2(n9465), .C1(n8197), .C2(n9462), .A(n1033), 
        .ZN(n1030) );
  AOI22_X1 U1435 ( .A1(n9459), .A2(n10113), .B1(n9454), .B2(n10145), .ZN(n1033) );
  OAI221_X1 U1436 ( .B1(n8316), .B2(n9465), .C1(n8187), .C2(n9462), .A(n943), 
        .ZN(n940) );
  AOI22_X1 U1437 ( .A1(n9459), .A2(n10108), .B1(n9454), .B2(n10140), .ZN(n943)
         );
  OAI221_X1 U1438 ( .B1(n8657), .B2(n9475), .C1(n8633), .C2(n9472), .A(n1410), 
        .ZN(n1409) );
  AOI22_X1 U1439 ( .A1(n9469), .A2(n10190), .B1(n9468), .B2(n10254), .ZN(n1410) );
  OAI221_X1 U1440 ( .B1(n8685), .B2(n9477), .C1(n8302), .C2(n9474), .A(n892), 
        .ZN(n889) );
  AOI22_X1 U1441 ( .A1(n9471), .A2(n10578), .B1(n9466), .B2(n10226), .ZN(n892)
         );
  OAI221_X1 U1442 ( .B1(n8668), .B2(n9476), .C1(n8644), .C2(n9473), .A(n1212), 
        .ZN(n1211) );
  AOI22_X1 U1443 ( .A1(n9470), .A2(n10179), .B1(n9467), .B2(n10243), .ZN(n1212) );
  OAI221_X1 U1444 ( .B1(n8664), .B2(n9475), .C1(n8640), .C2(n9472), .A(n1284), 
        .ZN(n1283) );
  AOI22_X1 U1445 ( .A1(n9469), .A2(n10183), .B1(n9467), .B2(n10247), .ZN(n1284) );
  OAI221_X1 U1446 ( .B1(n8672), .B2(n9476), .C1(n8648), .C2(n9473), .A(n1140), 
        .ZN(n1139) );
  AOI22_X1 U1447 ( .A1(n9470), .A2(n10175), .B1(n9467), .B2(n10239), .ZN(n1140) );
  OAI221_X1 U1448 ( .B1(n8682), .B2(n9477), .C1(n8299), .C2(n9474), .A(n960), 
        .ZN(n959) );
  AOI22_X1 U1449 ( .A1(n9471), .A2(n10581), .B1(n9466), .B2(n10229), .ZN(n960)
         );
  OAI221_X1 U1450 ( .B1(n8678), .B2(n9477), .C1(n8295), .C2(n9474), .A(n1032), 
        .ZN(n1031) );
  AOI22_X1 U1451 ( .A1(n9471), .A2(n10585), .B1(n9466), .B2(n10233), .ZN(n1032) );
  OAI221_X1 U1452 ( .B1(n8683), .B2(n9477), .C1(n8300), .C2(n9474), .A(n942), 
        .ZN(n941) );
  AOI22_X1 U1453 ( .A1(n9471), .A2(n10580), .B1(n9466), .B2(n10228), .ZN(n942)
         );
  AND3_X1 U1454 ( .A1(RD2), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n2077) );
  AND3_X1 U1455 ( .A1(RD2), .A2(n10661), .A3(ADD_RD2[3]), .ZN(n2095) );
  AND3_X1 U1456 ( .A1(n10662), .A2(n10661), .A3(RD2), .ZN(n2098) );
  OAI22_X1 U1457 ( .A1(n9870), .A2(n9259), .B1(n2157), .B2(n9867), .ZN(n9198)
         );
  OAI22_X1 U1458 ( .A1(n9870), .A2(n9256), .B1(n2149), .B2(n9868), .ZN(n9199)
         );
  OAI22_X1 U1459 ( .A1(n9870), .A2(n9253), .B1(n2141), .B2(n9867), .ZN(n9200)
         );
  OAI22_X1 U1460 ( .A1(n9869), .A2(n9250), .B1(n2133), .B2(n9868), .ZN(n9201)
         );
  OAI22_X1 U1461 ( .A1(n9869), .A2(n9247), .B1(n2125), .B2(n9867), .ZN(n9202)
         );
  OAI22_X1 U1462 ( .A1(n9869), .A2(n9244), .B1(n2117), .B2(n9868), .ZN(n9203)
         );
  OAI22_X1 U1463 ( .A1(n9869), .A2(n9241), .B1(n2109), .B2(n9867), .ZN(n9204)
         );
  OAI22_X1 U1464 ( .A1(n9869), .A2(n9238), .B1(n2101), .B2(n9868), .ZN(n9205)
         );
  OAI221_X1 U1465 ( .B1(n2327), .B2(n9487), .C1(n8378), .C2(n9484), .A(n1405), 
        .ZN(n1398) );
  AOI22_X1 U1466 ( .A1(n9481), .A2(n10222), .B1(n9480), .B2(n10654), .ZN(n1405) );
  AOI22_X1 U1467 ( .A1(n9505), .A2(n10606), .B1(n9504), .B2(n10438), .ZN(n1403) );
  OAI221_X1 U1468 ( .B1(n8629), .B2(n9525), .C1(n8597), .C2(n9522), .A(n868), 
        .ZN(n865) );
  AOI22_X1 U1469 ( .A1(n9519), .A2(n10442), .B1(n9514), .B2(n10258), .ZN(n868)
         );
  OAI221_X1 U1470 ( .B1(n2319), .B2(n9487), .C1(n8379), .C2(n9484), .A(n1387), 
        .ZN(n1380) );
  AOI22_X1 U1471 ( .A1(n9481), .A2(n10221), .B1(n9480), .B2(n10653), .ZN(n1387) );
  AOI22_X1 U1472 ( .A1(n9505), .A2(n10605), .B1(n9504), .B2(n10437), .ZN(n1385) );
  OAI221_X1 U1473 ( .B1(n2311), .B2(n9487), .C1(n8380), .C2(n9484), .A(n1369), 
        .ZN(n1362) );
  AOI22_X1 U1474 ( .A1(n9481), .A2(n10220), .B1(n9480), .B2(n10652), .ZN(n1369) );
  AOI22_X1 U1475 ( .A1(n9505), .A2(n10604), .B1(n9504), .B2(n10436), .ZN(n1367) );
  OAI221_X1 U1476 ( .B1(n8611), .B2(n9524), .C1(n8579), .C2(n9521), .A(n1222), 
        .ZN(n1221) );
  AOI22_X1 U1477 ( .A1(n9518), .A2(n10460), .B1(n9515), .B2(n10276), .ZN(n1222) );
  OAI221_X1 U1478 ( .B1(n8612), .B2(n9524), .C1(n8580), .C2(n9521), .A(n1204), 
        .ZN(n1203) );
  AOI22_X1 U1479 ( .A1(n9518), .A2(n10459), .B1(n9515), .B2(n10275), .ZN(n1204) );
  OAI221_X1 U1480 ( .B1(n8613), .B2(n9524), .C1(n8581), .C2(n9521), .A(n1186), 
        .ZN(n1185) );
  AOI22_X1 U1481 ( .A1(n9518), .A2(n10458), .B1(n9515), .B2(n10274), .ZN(n1186) );
  OAI221_X1 U1482 ( .B1(n2351), .B2(n9487), .C1(n8375), .C2(n9484), .A(n1469), 
        .ZN(n1452) );
  AOI22_X1 U1483 ( .A1(n9481), .A2(n10225), .B1(n9480), .B2(n10657), .ZN(n1469) );
  OAI221_X1 U1484 ( .B1(n8252), .B2(n9512), .C1(n8218), .C2(n9509), .A(n1223), 
        .ZN(n1220) );
  AOI22_X1 U1485 ( .A1(n9506), .A2(n10596), .B1(n9503), .B2(n10428), .ZN(n1223) );
  AOI22_X1 U1486 ( .A1(n9434), .A2(n10332), .B1(n9431), .B2(n9940), .ZN(n1233)
         );
  AOI22_X1 U1487 ( .A1(n9433), .A2(n10345), .B1(n9432), .B2(n9953), .ZN(n1479)
         );
  AOI22_X1 U1488 ( .A1(n9506), .A2(n10595), .B1(n9503), .B2(n10427), .ZN(n1205) );
  AOI22_X1 U1489 ( .A1(n9506), .A2(n10594), .B1(n9503), .B2(n10426), .ZN(n1187) );
  AOI22_X1 U1490 ( .A1(n9506), .A2(n10589), .B1(n9502), .B2(n10421), .ZN(n1097) );
  AOI22_X1 U1491 ( .A1(n9505), .A2(n10599), .B1(n9503), .B2(n10431), .ZN(n1277) );
  AOI22_X1 U1492 ( .A1(n9505), .A2(n10598), .B1(n9503), .B2(n10430), .ZN(n1259) );
  AOI22_X1 U1493 ( .A1(n9506), .A2(n10587), .B1(n9502), .B2(n10419), .ZN(n1061) );
  AOI22_X1 U1494 ( .A1(n9506), .A2(n10588), .B1(n9502), .B2(n10420), .ZN(n1079) );
  AOI22_X1 U1495 ( .A1(n9506), .A2(n10593), .B1(n9503), .B2(n10425), .ZN(n1169) );
  AOI22_X1 U1496 ( .A1(n9506), .A2(n10597), .B1(n9503), .B2(n10429), .ZN(n1241) );
  AOI22_X1 U1497 ( .A1(n9506), .A2(n10586), .B1(n9502), .B2(n10418), .ZN(n1043) );
  OAI221_X1 U1498 ( .B1(n8615), .B2(n9524), .C1(n8583), .C2(n9521), .A(n1150), 
        .ZN(n1149) );
  AOI22_X1 U1499 ( .A1(n9518), .A2(n10456), .B1(n9515), .B2(n10272), .ZN(n1150) );
  OAI221_X1 U1500 ( .B1(n8616), .B2(n9524), .C1(n8584), .C2(n9521), .A(n1132), 
        .ZN(n1131) );
  AOI22_X1 U1501 ( .A1(n9518), .A2(n10455), .B1(n9515), .B2(n10271), .ZN(n1132) );
  OAI221_X1 U1502 ( .B1(n8617), .B2(n9524), .C1(n8585), .C2(n9521), .A(n1114), 
        .ZN(n1113) );
  AOI22_X1 U1503 ( .A1(n9518), .A2(n10454), .B1(n9515), .B2(n10270), .ZN(n1114) );
  OAI221_X1 U1504 ( .B1(n8256), .B2(n9512), .C1(n8210), .C2(n9509), .A(n1151), 
        .ZN(n1148) );
  AOI22_X1 U1505 ( .A1(n9506), .A2(n10592), .B1(n9503), .B2(n10424), .ZN(n1151) );
  AOI22_X1 U1506 ( .A1(n9434), .A2(n10328), .B1(n9431), .B2(n9936), .ZN(n1161)
         );
  AOI22_X1 U1507 ( .A1(n9506), .A2(n10591), .B1(n9503), .B2(n10423), .ZN(n1133) );
  AOI22_X1 U1508 ( .A1(n9506), .A2(n10590), .B1(n9503), .B2(n10422), .ZN(n1115) );
  OAI221_X1 U1509 ( .B1(n2343), .B2(n9487), .C1(n8376), .C2(n9484), .A(n1441), 
        .ZN(n1434) );
  AOI22_X1 U1510 ( .A1(n9481), .A2(n10224), .B1(n9480), .B2(n10656), .ZN(n1441) );
  AOI22_X1 U1511 ( .A1(n9505), .A2(n10608), .B1(n9504), .B2(n10440), .ZN(n1439) );
  OAI221_X1 U1512 ( .B1(n8623), .B2(n9525), .C1(n8591), .C2(n9522), .A(n1006), 
        .ZN(n1005) );
  AOI22_X1 U1513 ( .A1(n9519), .A2(n10448), .B1(n9514), .B2(n10264), .ZN(n1006) );
  OAI221_X1 U1514 ( .B1(n8626), .B2(n9525), .C1(n8594), .C2(n9522), .A(n952), 
        .ZN(n951) );
  AOI22_X1 U1515 ( .A1(n9519), .A2(n10445), .B1(n9514), .B2(n10261), .ZN(n952)
         );
  OAI221_X1 U1516 ( .B1(n2335), .B2(n9487), .C1(n8377), .C2(n9484), .A(n1423), 
        .ZN(n1416) );
  AOI22_X1 U1517 ( .A1(n9481), .A2(n10223), .B1(n9480), .B2(n10655), .ZN(n1423) );
  OAI221_X1 U1518 ( .B1(n2303), .B2(n9487), .C1(n8381), .C2(n9484), .A(n1351), 
        .ZN(n1344) );
  AOI22_X1 U1519 ( .A1(n9481), .A2(n10219), .B1(n9480), .B2(n10651), .ZN(n1351) );
  OAI221_X1 U1520 ( .B1(n2295), .B2(n9487), .C1(n8382), .C2(n9484), .A(n1333), 
        .ZN(n1326) );
  AOI22_X1 U1521 ( .A1(n9481), .A2(n10218), .B1(n9480), .B2(n10650), .ZN(n1333) );
  AOI22_X1 U1522 ( .A1(n9505), .A2(n10607), .B1(n9504), .B2(n10439), .ZN(n1421) );
  AOI22_X1 U1523 ( .A1(n9433), .A2(n10339), .B1(n9432), .B2(n9947), .ZN(n1359)
         );
  AOI22_X1 U1524 ( .A1(n9505), .A2(n10602), .B1(n9504), .B2(n10434), .ZN(n1331) );
  AOI22_X1 U1525 ( .A1(n9505), .A2(n10601), .B1(n9503), .B2(n10433), .ZN(n1313) );
  AOI22_X1 U1526 ( .A1(n9505), .A2(n10600), .B1(n9503), .B2(n10432), .ZN(n1295) );
  AOI22_X1 U1527 ( .A1(n9349), .A2(n10041), .B1(n9348), .B2(n10073), .ZN(n2097) );
  AOI22_X1 U1528 ( .A1(n9361), .A2(n10105), .B1(n9360), .B2(n10137), .ZN(n2096) );
  AOI22_X1 U1529 ( .A1(n9337), .A2(n9953), .B1(n9336), .B2(n9985), .ZN(n2099)
         );
  AOI22_X1 U1530 ( .A1(n9349), .A2(n10040), .B1(n9348), .B2(n10072), .ZN(n2068) );
  AOI22_X1 U1531 ( .A1(n9361), .A2(n10104), .B1(n9360), .B2(n10136), .ZN(n2067) );
  AOI22_X1 U1532 ( .A1(n9337), .A2(n9952), .B1(n9336), .B2(n9984), .ZN(n2069)
         );
  AOI22_X1 U1533 ( .A1(n9349), .A2(n10039), .B1(n9348), .B2(n10071), .ZN(n2050) );
  AOI22_X1 U1534 ( .A1(n9361), .A2(n10103), .B1(n9360), .B2(n10135), .ZN(n2049) );
  AOI22_X1 U1535 ( .A1(n9337), .A2(n9951), .B1(n9336), .B2(n9983), .ZN(n2051)
         );
  AOI22_X1 U1536 ( .A1(n9349), .A2(n10038), .B1(n9348), .B2(n10070), .ZN(n2032) );
  AOI22_X1 U1537 ( .A1(n9361), .A2(n10102), .B1(n9360), .B2(n10134), .ZN(n2031) );
  AOI22_X1 U1538 ( .A1(n9337), .A2(n9950), .B1(n9336), .B2(n9982), .ZN(n2033)
         );
  AOI22_X1 U1539 ( .A1(n9349), .A2(n10037), .B1(n9348), .B2(n10069), .ZN(n2014) );
  AOI22_X1 U1540 ( .A1(n9361), .A2(n10101), .B1(n9360), .B2(n10133), .ZN(n2013) );
  AOI22_X1 U1541 ( .A1(n9337), .A2(n9949), .B1(n9336), .B2(n9981), .ZN(n2015)
         );
  AOI22_X1 U1542 ( .A1(n9349), .A2(n10036), .B1(n9348), .B2(n10068), .ZN(n1996) );
  AOI22_X1 U1543 ( .A1(n9361), .A2(n10100), .B1(n9360), .B2(n10132), .ZN(n1995) );
  AOI22_X1 U1544 ( .A1(n9337), .A2(n9948), .B1(n9336), .B2(n9980), .ZN(n1997)
         );
  AOI22_X1 U1545 ( .A1(n9349), .A2(n10035), .B1(n9348), .B2(n10067), .ZN(n1978) );
  AOI22_X1 U1546 ( .A1(n9361), .A2(n10099), .B1(n9360), .B2(n10131), .ZN(n1977) );
  AOI22_X1 U1547 ( .A1(n9337), .A2(n9947), .B1(n9336), .B2(n9979), .ZN(n1979)
         );
  AOI22_X1 U1548 ( .A1(n9349), .A2(n10034), .B1(n9348), .B2(n10066), .ZN(n1960) );
  AOI22_X1 U1549 ( .A1(n9361), .A2(n10098), .B1(n9360), .B2(n10130), .ZN(n1959) );
  AOI22_X1 U1550 ( .A1(n9337), .A2(n9946), .B1(n9336), .B2(n9978), .ZN(n1961)
         );
  AOI22_X1 U1551 ( .A1(n9409), .A2(n10625), .B1(n9407), .B2(n10601), .ZN(n1933) );
  AOI22_X1 U1552 ( .A1(n9397), .A2(n10369), .B1(n9395), .B2(n10401), .ZN(n1934) );
  AOI22_X1 U1553 ( .A1(n9385), .A2(n10281), .B1(n9383), .B2(n10313), .ZN(n1935) );
  AOI22_X1 U1554 ( .A1(n9409), .A2(n10624), .B1(n9407), .B2(n10600), .ZN(n1915) );
  AOI22_X1 U1555 ( .A1(n9397), .A2(n10368), .B1(n9395), .B2(n10400), .ZN(n1916) );
  AOI22_X1 U1556 ( .A1(n9385), .A2(n10280), .B1(n9383), .B2(n10312), .ZN(n1917) );
  AOI22_X1 U1557 ( .A1(n9409), .A2(n10623), .B1(n9407), .B2(n10599), .ZN(n1897) );
  AOI22_X1 U1558 ( .A1(n9397), .A2(n10367), .B1(n9395), .B2(n10399), .ZN(n1898) );
  AOI22_X1 U1559 ( .A1(n9385), .A2(n10279), .B1(n9383), .B2(n10311), .ZN(n1899) );
  AOI22_X1 U1560 ( .A1(n9409), .A2(n10622), .B1(n9407), .B2(n10598), .ZN(n1879) );
  AOI22_X1 U1561 ( .A1(n9397), .A2(n10366), .B1(n9395), .B2(n10398), .ZN(n1880) );
  AOI22_X1 U1562 ( .A1(n9385), .A2(n10278), .B1(n9383), .B2(n10310), .ZN(n1881) );
  AOI22_X1 U1563 ( .A1(n9410), .A2(n10621), .B1(n9407), .B2(n10597), .ZN(n1861) );
  AOI22_X1 U1564 ( .A1(n9398), .A2(n10365), .B1(n9395), .B2(n10397), .ZN(n1862) );
  AOI22_X1 U1565 ( .A1(n9386), .A2(n10277), .B1(n9383), .B2(n10309), .ZN(n1863) );
  AOI22_X1 U1566 ( .A1(n9410), .A2(n10620), .B1(n9407), .B2(n10596), .ZN(n1843) );
  AOI22_X1 U1567 ( .A1(n9398), .A2(n10364), .B1(n9395), .B2(n10396), .ZN(n1844) );
  AOI22_X1 U1568 ( .A1(n9386), .A2(n10276), .B1(n9383), .B2(n10308), .ZN(n1845) );
  AOI22_X1 U1569 ( .A1(n9410), .A2(n10619), .B1(n9407), .B2(n10595), .ZN(n1825) );
  AOI22_X1 U1570 ( .A1(n9398), .A2(n10363), .B1(n9395), .B2(n10395), .ZN(n1826) );
  AOI22_X1 U1571 ( .A1(n9386), .A2(n10275), .B1(n9383), .B2(n10307), .ZN(n1827) );
  AOI22_X1 U1572 ( .A1(n9410), .A2(n10618), .B1(n9407), .B2(n10594), .ZN(n1807) );
  AOI22_X1 U1573 ( .A1(n9398), .A2(n10362), .B1(n9395), .B2(n10394), .ZN(n1808) );
  AOI22_X1 U1574 ( .A1(n9386), .A2(n10274), .B1(n9383), .B2(n10306), .ZN(n1809) );
  AOI22_X1 U1575 ( .A1(n9410), .A2(n10617), .B1(n9407), .B2(n10593), .ZN(n1789) );
  AOI22_X1 U1576 ( .A1(n9398), .A2(n10361), .B1(n9395), .B2(n10393), .ZN(n1790) );
  AOI22_X1 U1577 ( .A1(n9386), .A2(n10273), .B1(n9383), .B2(n10305), .ZN(n1791) );
  AOI22_X1 U1578 ( .A1(n9410), .A2(n10616), .B1(n9407), .B2(n10592), .ZN(n1771) );
  AOI22_X1 U1579 ( .A1(n9398), .A2(n10360), .B1(n9395), .B2(n10392), .ZN(n1772) );
  AOI22_X1 U1580 ( .A1(n9386), .A2(n10272), .B1(n9383), .B2(n10304), .ZN(n1773) );
  AOI22_X1 U1581 ( .A1(n9410), .A2(n10615), .B1(n9407), .B2(n10591), .ZN(n1753) );
  AOI22_X1 U1582 ( .A1(n9398), .A2(n10359), .B1(n9395), .B2(n10391), .ZN(n1754) );
  AOI22_X1 U1583 ( .A1(n9386), .A2(n10271), .B1(n9383), .B2(n10303), .ZN(n1755) );
  AOI22_X1 U1584 ( .A1(n9410), .A2(n10614), .B1(n9407), .B2(n10590), .ZN(n1735) );
  AOI22_X1 U1585 ( .A1(n9398), .A2(n10358), .B1(n9395), .B2(n10390), .ZN(n1736) );
  AOI22_X1 U1586 ( .A1(n9386), .A2(n10270), .B1(n9383), .B2(n10302), .ZN(n1737) );
  AOI22_X1 U1587 ( .A1(n9410), .A2(n10613), .B1(n9406), .B2(n10589), .ZN(n1717) );
  AOI22_X1 U1588 ( .A1(n9398), .A2(n10357), .B1(n9394), .B2(n10389), .ZN(n1718) );
  AOI22_X1 U1589 ( .A1(n9386), .A2(n10269), .B1(n9382), .B2(n10301), .ZN(n1719) );
  AOI22_X1 U1590 ( .A1(n9410), .A2(n10612), .B1(n9406), .B2(n10588), .ZN(n1699) );
  AOI22_X1 U1591 ( .A1(n9398), .A2(n10356), .B1(n9394), .B2(n10388), .ZN(n1700) );
  AOI22_X1 U1592 ( .A1(n9386), .A2(n10268), .B1(n9382), .B2(n10300), .ZN(n1701) );
  AOI22_X1 U1593 ( .A1(n9410), .A2(n10611), .B1(n9406), .B2(n10587), .ZN(n1681) );
  AOI22_X1 U1594 ( .A1(n9398), .A2(n10355), .B1(n9394), .B2(n10387), .ZN(n1682) );
  AOI22_X1 U1595 ( .A1(n9386), .A2(n10267), .B1(n9382), .B2(n10299), .ZN(n1683) );
  AOI22_X1 U1596 ( .A1(n9410), .A2(n10610), .B1(n9406), .B2(n10586), .ZN(n1663) );
  AOI22_X1 U1597 ( .A1(n9398), .A2(n10354), .B1(n9394), .B2(n10386), .ZN(n1664) );
  AOI22_X1 U1598 ( .A1(n9386), .A2(n10266), .B1(n9382), .B2(n10298), .ZN(n1665) );
  AOI22_X1 U1599 ( .A1(n9411), .A2(n10553), .B1(n9406), .B2(n10545), .ZN(n1645) );
  AOI22_X1 U1600 ( .A1(n9399), .A2(n10353), .B1(n9394), .B2(n10385), .ZN(n1646) );
  AOI22_X1 U1601 ( .A1(n9387), .A2(n10265), .B1(n9382), .B2(n10297), .ZN(n1647) );
  AOI22_X1 U1602 ( .A1(n9411), .A2(n10552), .B1(n9406), .B2(n10544), .ZN(n1627) );
  AOI22_X1 U1603 ( .A1(n9399), .A2(n10352), .B1(n9394), .B2(n10384), .ZN(n1628) );
  AOI22_X1 U1604 ( .A1(n9387), .A2(n10264), .B1(n9382), .B2(n10296), .ZN(n1629) );
  AOI22_X1 U1605 ( .A1(n9411), .A2(n10551), .B1(n9406), .B2(n10543), .ZN(n1609) );
  AOI22_X1 U1606 ( .A1(n9399), .A2(n10351), .B1(n9394), .B2(n10383), .ZN(n1610) );
  AOI22_X1 U1607 ( .A1(n9387), .A2(n10263), .B1(n9382), .B2(n10295), .ZN(n1611) );
  AOI22_X1 U1608 ( .A1(n9411), .A2(n10550), .B1(n9406), .B2(n10542), .ZN(n1591) );
  AOI22_X1 U1609 ( .A1(n9399), .A2(n10350), .B1(n9394), .B2(n10382), .ZN(n1592) );
  AOI22_X1 U1610 ( .A1(n9387), .A2(n10262), .B1(n9382), .B2(n10294), .ZN(n1593) );
  AOI22_X1 U1611 ( .A1(n9411), .A2(n10549), .B1(n9406), .B2(n10541), .ZN(n1573) );
  AOI22_X1 U1612 ( .A1(n9399), .A2(n10349), .B1(n9394), .B2(n10381), .ZN(n1574) );
  AOI22_X1 U1613 ( .A1(n9387), .A2(n10261), .B1(n9382), .B2(n10293), .ZN(n1575) );
  AOI22_X1 U1614 ( .A1(n9411), .A2(n10548), .B1(n9406), .B2(n10540), .ZN(n1555) );
  AOI22_X1 U1615 ( .A1(n9399), .A2(n10348), .B1(n9394), .B2(n10380), .ZN(n1556) );
  AOI22_X1 U1616 ( .A1(n9387), .A2(n10260), .B1(n9382), .B2(n10292), .ZN(n1557) );
  AOI22_X1 U1617 ( .A1(n9411), .A2(n10547), .B1(n9406), .B2(n10539), .ZN(n1537) );
  AOI22_X1 U1618 ( .A1(n9399), .A2(n10347), .B1(n9394), .B2(n10379), .ZN(n1538) );
  AOI22_X1 U1619 ( .A1(n9387), .A2(n10259), .B1(n9382), .B2(n10291), .ZN(n1539) );
  AOI22_X1 U1620 ( .A1(n9411), .A2(n10546), .B1(n9406), .B2(n10538), .ZN(n1493) );
  AOI22_X1 U1621 ( .A1(n9399), .A2(n10346), .B1(n9394), .B2(n10378), .ZN(n1498) );
  AOI22_X1 U1622 ( .A1(n9387), .A2(n10258), .B1(n9382), .B2(n10290), .ZN(n1503) );
  OAI221_X1 U1623 ( .B1(n8654), .B2(n9379), .C1(n8630), .C2(n9376), .A(n2094), 
        .ZN(n2093) );
  AOI22_X1 U1624 ( .A1(n9373), .A2(n10225), .B1(n9372), .B2(n10257), .ZN(n2094) );
  OAI221_X1 U1625 ( .B1(n8375), .B2(n9427), .C1(n8343), .C2(n9424), .A(n2076), 
        .ZN(n2075) );
  AOI22_X1 U1626 ( .A1(n9421), .A2(n10657), .B1(n9420), .B2(n10537), .ZN(n2076) );
  OAI221_X1 U1627 ( .B1(n8439), .B2(n9415), .C1(n8407), .C2(n9412), .A(n2082), 
        .ZN(n2074) );
  AOI22_X1 U1628 ( .A1(n9409), .A2(n10633), .B1(n9408), .B2(n10609), .ZN(n2082) );
  OAI221_X1 U1629 ( .B1(n8478), .B2(n9403), .C1(n8471), .C2(n9400), .A(n2087), 
        .ZN(n2073) );
  AOI22_X1 U1630 ( .A1(n9397), .A2(n10377), .B1(n9396), .B2(n10409), .ZN(n2087) );
  OAI221_X1 U1631 ( .B1(n8566), .B2(n9391), .C1(n8542), .C2(n9388), .A(n2089), 
        .ZN(n2072) );
  AOI22_X1 U1632 ( .A1(n9385), .A2(n10289), .B1(n9384), .B2(n10321), .ZN(n2089) );
  OAI221_X1 U1633 ( .B1(n8655), .B2(n9379), .C1(n8631), .C2(n9376), .A(n2066), 
        .ZN(n2065) );
  AOI22_X1 U1634 ( .A1(n9373), .A2(n10224), .B1(n9372), .B2(n10256), .ZN(n2066) );
  OAI221_X1 U1635 ( .B1(n8376), .B2(n9427), .C1(n8344), .C2(n9424), .A(n2058), 
        .ZN(n2057) );
  AOI22_X1 U1636 ( .A1(n9421), .A2(n10656), .B1(n9420), .B2(n10536), .ZN(n2058) );
  OAI221_X1 U1637 ( .B1(n8440), .B2(n9415), .C1(n8408), .C2(n9412), .A(n2059), 
        .ZN(n2056) );
  AOI22_X1 U1638 ( .A1(n9409), .A2(n10632), .B1(n9408), .B2(n10608), .ZN(n2059) );
  OAI221_X1 U1639 ( .B1(n8479), .B2(n9403), .C1(n8472), .C2(n9400), .A(n2060), 
        .ZN(n2055) );
  AOI22_X1 U1640 ( .A1(n9397), .A2(n10376), .B1(n9396), .B2(n10408), .ZN(n2060) );
  OAI221_X1 U1641 ( .B1(n8567), .B2(n9391), .C1(n8543), .C2(n9388), .A(n2061), 
        .ZN(n2054) );
  AOI22_X1 U1642 ( .A1(n9385), .A2(n10288), .B1(n9384), .B2(n10320), .ZN(n2061) );
  OAI221_X1 U1643 ( .B1(n8656), .B2(n9379), .C1(n8632), .C2(n9376), .A(n2048), 
        .ZN(n2047) );
  AOI22_X1 U1644 ( .A1(n9373), .A2(n10223), .B1(n9372), .B2(n10255), .ZN(n2048) );
  OAI221_X1 U1645 ( .B1(n8377), .B2(n9427), .C1(n8345), .C2(n9424), .A(n2040), 
        .ZN(n2039) );
  AOI22_X1 U1646 ( .A1(n9421), .A2(n10655), .B1(n9420), .B2(n10535), .ZN(n2040) );
  OAI221_X1 U1647 ( .B1(n8441), .B2(n9415), .C1(n8409), .C2(n9412), .A(n2041), 
        .ZN(n2038) );
  AOI22_X1 U1648 ( .A1(n9409), .A2(n10631), .B1(n9408), .B2(n10607), .ZN(n2041) );
  OAI221_X1 U1649 ( .B1(n8480), .B2(n9403), .C1(n8473), .C2(n9400), .A(n2042), 
        .ZN(n2037) );
  AOI22_X1 U1650 ( .A1(n9397), .A2(n10375), .B1(n9396), .B2(n10407), .ZN(n2042) );
  OAI221_X1 U1651 ( .B1(n8568), .B2(n9391), .C1(n8544), .C2(n9388), .A(n2043), 
        .ZN(n2036) );
  AOI22_X1 U1652 ( .A1(n9385), .A2(n10287), .B1(n9384), .B2(n10319), .ZN(n2043) );
  OAI221_X1 U1653 ( .B1(n8657), .B2(n9379), .C1(n8633), .C2(n9376), .A(n2030), 
        .ZN(n2029) );
  AOI22_X1 U1654 ( .A1(n9373), .A2(n10222), .B1(n9372), .B2(n10254), .ZN(n2030) );
  OAI221_X1 U1655 ( .B1(n8378), .B2(n9427), .C1(n8346), .C2(n9424), .A(n2022), 
        .ZN(n2021) );
  AOI22_X1 U1656 ( .A1(n9421), .A2(n10654), .B1(n9420), .B2(n10534), .ZN(n2022) );
  OAI221_X1 U1657 ( .B1(n8442), .B2(n9415), .C1(n8410), .C2(n9412), .A(n2023), 
        .ZN(n2020) );
  AOI22_X1 U1658 ( .A1(n9409), .A2(n10630), .B1(n9408), .B2(n10606), .ZN(n2023) );
  OAI221_X1 U1659 ( .B1(n8481), .B2(n9403), .C1(n8474), .C2(n9400), .A(n2024), 
        .ZN(n2019) );
  AOI22_X1 U1660 ( .A1(n9397), .A2(n10374), .B1(n9396), .B2(n10406), .ZN(n2024) );
  OAI221_X1 U1661 ( .B1(n8569), .B2(n9391), .C1(n8545), .C2(n9388), .A(n2025), 
        .ZN(n2018) );
  AOI22_X1 U1662 ( .A1(n9385), .A2(n10286), .B1(n9384), .B2(n10318), .ZN(n2025) );
  OAI221_X1 U1663 ( .B1(n8658), .B2(n9379), .C1(n8634), .C2(n9376), .A(n2012), 
        .ZN(n2011) );
  AOI22_X1 U1664 ( .A1(n9373), .A2(n10221), .B1(n9372), .B2(n10253), .ZN(n2012) );
  OAI221_X1 U1665 ( .B1(n8379), .B2(n9427), .C1(n8347), .C2(n9424), .A(n2004), 
        .ZN(n2003) );
  AOI22_X1 U1666 ( .A1(n9421), .A2(n10653), .B1(n9420), .B2(n10533), .ZN(n2004) );
  OAI221_X1 U1667 ( .B1(n8443), .B2(n9415), .C1(n8411), .C2(n9412), .A(n2005), 
        .ZN(n2002) );
  AOI22_X1 U1668 ( .A1(n9409), .A2(n10629), .B1(n9408), .B2(n10605), .ZN(n2005) );
  OAI221_X1 U1669 ( .B1(n8482), .B2(n9403), .C1(n8475), .C2(n9400), .A(n2006), 
        .ZN(n2001) );
  AOI22_X1 U1670 ( .A1(n9397), .A2(n10373), .B1(n9396), .B2(n10405), .ZN(n2006) );
  OAI221_X1 U1671 ( .B1(n8570), .B2(n9391), .C1(n8546), .C2(n9388), .A(n2007), 
        .ZN(n2000) );
  AOI22_X1 U1672 ( .A1(n9385), .A2(n10285), .B1(n9384), .B2(n10317), .ZN(n2007) );
  OAI221_X1 U1673 ( .B1(n8659), .B2(n9379), .C1(n8635), .C2(n9376), .A(n1994), 
        .ZN(n1993) );
  AOI22_X1 U1674 ( .A1(n9373), .A2(n10220), .B1(n9372), .B2(n10252), .ZN(n1994) );
  OAI221_X1 U1675 ( .B1(n8380), .B2(n9427), .C1(n8348), .C2(n9424), .A(n1986), 
        .ZN(n1985) );
  AOI22_X1 U1676 ( .A1(n9421), .A2(n10652), .B1(n9420), .B2(n10532), .ZN(n1986) );
  OAI221_X1 U1677 ( .B1(n8444), .B2(n9415), .C1(n8412), .C2(n9412), .A(n1987), 
        .ZN(n1984) );
  AOI22_X1 U1678 ( .A1(n9409), .A2(n10628), .B1(n9408), .B2(n10604), .ZN(n1987) );
  OAI221_X1 U1679 ( .B1(n8483), .B2(n9403), .C1(n8476), .C2(n9400), .A(n1988), 
        .ZN(n1983) );
  AOI22_X1 U1680 ( .A1(n9397), .A2(n10372), .B1(n9396), .B2(n10404), .ZN(n1988) );
  OAI221_X1 U1681 ( .B1(n8571), .B2(n9391), .C1(n8547), .C2(n9388), .A(n1989), 
        .ZN(n1982) );
  AOI22_X1 U1682 ( .A1(n9385), .A2(n10284), .B1(n9384), .B2(n10316), .ZN(n1989) );
  OAI221_X1 U1683 ( .B1(n8660), .B2(n9379), .C1(n8636), .C2(n9376), .A(n1976), 
        .ZN(n1975) );
  AOI22_X1 U1684 ( .A1(n9373), .A2(n10219), .B1(n9372), .B2(n10251), .ZN(n1976) );
  OAI221_X1 U1685 ( .B1(n8381), .B2(n9427), .C1(n8349), .C2(n9424), .A(n1968), 
        .ZN(n1967) );
  AOI22_X1 U1687 ( .A1(n9421), .A2(n10651), .B1(n9420), .B2(n10531), .ZN(n1968) );
  OAI221_X1 U1688 ( .B1(n8445), .B2(n9415), .C1(n8413), .C2(n9412), .A(n1969), 
        .ZN(n1966) );
  AOI22_X1 U1689 ( .A1(n9409), .A2(n10627), .B1(n9408), .B2(n10603), .ZN(n1969) );
  OAI221_X1 U1690 ( .B1(n8484), .B2(n9403), .C1(n8477), .C2(n9400), .A(n1970), 
        .ZN(n1965) );
  AOI22_X1 U1691 ( .A1(n9397), .A2(n10371), .B1(n9396), .B2(n10403), .ZN(n1970) );
  OAI221_X1 U1692 ( .B1(n8572), .B2(n9391), .C1(n8548), .C2(n9388), .A(n1971), 
        .ZN(n1964) );
  AOI22_X1 U1693 ( .A1(n9385), .A2(n10283), .B1(n9384), .B2(n10315), .ZN(n1971) );
  OAI221_X1 U1694 ( .B1(n8661), .B2(n9379), .C1(n8637), .C2(n9376), .A(n1958), 
        .ZN(n1957) );
  AOI22_X1 U1695 ( .A1(n9373), .A2(n10218), .B1(n9372), .B2(n10250), .ZN(n1958) );
  OAI221_X1 U1696 ( .B1(n8382), .B2(n9427), .C1(n8350), .C2(n9424), .A(n1950), 
        .ZN(n1949) );
  AOI22_X1 U1697 ( .A1(n9421), .A2(n10650), .B1(n9420), .B2(n10530), .ZN(n1950) );
  OAI221_X1 U1698 ( .B1(n8446), .B2(n9415), .C1(n8414), .C2(n9412), .A(n1951), 
        .ZN(n1948) );
  AOI22_X1 U1700 ( .A1(n9409), .A2(n10626), .B1(n9408), .B2(n10602), .ZN(n1951) );
  OAI221_X1 U1701 ( .B1(n8485), .B2(n9403), .C1(n8246), .C2(n9400), .A(n1952), 
        .ZN(n1947) );
  AOI22_X1 U1702 ( .A1(n9397), .A2(n10370), .B1(n9396), .B2(n10402), .ZN(n1952) );
  OAI221_X1 U1703 ( .B1(n8573), .B2(n9391), .C1(n8549), .C2(n9388), .A(n1953), 
        .ZN(n1946) );
  AOI22_X1 U1704 ( .A1(n9385), .A2(n10282), .B1(n9384), .B2(n10314), .ZN(n1953) );
  OAI221_X1 U1705 ( .B1(n8383), .B2(n9427), .C1(n8351), .C2(n9424), .A(n1932), 
        .ZN(n1931) );
  AOI22_X1 U1706 ( .A1(n9421), .A2(n10649), .B1(n9419), .B2(n10529), .ZN(n1932) );
  OAI221_X1 U1707 ( .B1(n8750), .B2(n9367), .C1(n8726), .C2(n9364), .A(n1941), 
        .ZN(n1938) );
  AOI22_X1 U1708 ( .A1(n9361), .A2(n10097), .B1(n9359), .B2(n10129), .ZN(n1941) );
  OAI221_X1 U1709 ( .B1(n8384), .B2(n9427), .C1(n8352), .C2(n9424), .A(n1914), 
        .ZN(n1913) );
  AOI22_X1 U1710 ( .A1(n9421), .A2(n10648), .B1(n9419), .B2(n10528), .ZN(n1914) );
  OAI221_X1 U1711 ( .B1(n8751), .B2(n9367), .C1(n8727), .C2(n9364), .A(n1923), 
        .ZN(n1920) );
  AOI22_X1 U1712 ( .A1(n9361), .A2(n10096), .B1(n9359), .B2(n10128), .ZN(n1923) );
  OAI221_X1 U1713 ( .B1(n8385), .B2(n9427), .C1(n8353), .C2(n9424), .A(n1896), 
        .ZN(n1895) );
  AOI22_X1 U1714 ( .A1(n9421), .A2(n10647), .B1(n9419), .B2(n10527), .ZN(n1896) );
  OAI221_X1 U1715 ( .B1(n8752), .B2(n9367), .C1(n8728), .C2(n9364), .A(n1905), 
        .ZN(n1902) );
  AOI22_X1 U1717 ( .A1(n9361), .A2(n10095), .B1(n9359), .B2(n10127), .ZN(n1905) );
  OAI221_X1 U1718 ( .B1(n8386), .B2(n9427), .C1(n8354), .C2(n9424), .A(n1878), 
        .ZN(n1877) );
  AOI22_X1 U1719 ( .A1(n9421), .A2(n10646), .B1(n9419), .B2(n10526), .ZN(n1878) );
  OAI221_X1 U1720 ( .B1(n8753), .B2(n9367), .C1(n8729), .C2(n9364), .A(n1887), 
        .ZN(n1884) );
  AOI22_X1 U1721 ( .A1(n9361), .A2(n10094), .B1(n9359), .B2(n10126), .ZN(n1887) );
  OAI221_X1 U1723 ( .B1(n8387), .B2(n9428), .C1(n8355), .C2(n9425), .A(n1860), 
        .ZN(n1859) );
  AOI22_X1 U1724 ( .A1(n9422), .A2(n10645), .B1(n9419), .B2(n10525), .ZN(n1860) );
  OAI221_X1 U1725 ( .B1(n8754), .B2(n9368), .C1(n8730), .C2(n9365), .A(n1869), 
        .ZN(n1866) );
  AOI22_X1 U1726 ( .A1(n9362), .A2(n10093), .B1(n9359), .B2(n10125), .ZN(n1869) );
  OAI221_X1 U1727 ( .B1(n8388), .B2(n9428), .C1(n8356), .C2(n9425), .A(n1842), 
        .ZN(n1841) );
  AOI22_X1 U1728 ( .A1(n9422), .A2(n10644), .B1(n9419), .B2(n10524), .ZN(n1842) );
  OAI221_X1 U1729 ( .B1(n8755), .B2(n9368), .C1(n8731), .C2(n9365), .A(n1851), 
        .ZN(n1848) );
  AOI22_X1 U1730 ( .A1(n9362), .A2(n10092), .B1(n9359), .B2(n10124), .ZN(n1851) );
  OAI221_X1 U1731 ( .B1(n8389), .B2(n9428), .C1(n8357), .C2(n9425), .A(n1824), 
        .ZN(n1823) );
  AOI22_X1 U1732 ( .A1(n9422), .A2(n10643), .B1(n9419), .B2(n10523), .ZN(n1824) );
  OAI221_X1 U1733 ( .B1(n8756), .B2(n9368), .C1(n8732), .C2(n9365), .A(n1833), 
        .ZN(n1830) );
  AOI22_X1 U1734 ( .A1(n9362), .A2(n10091), .B1(n9359), .B2(n10123), .ZN(n1833) );
  OAI221_X1 U1735 ( .B1(n8390), .B2(n9428), .C1(n8358), .C2(n9425), .A(n1806), 
        .ZN(n1805) );
  AOI22_X1 U1736 ( .A1(n9422), .A2(n10642), .B1(n9419), .B2(n10522), .ZN(n1806) );
  OAI221_X1 U1737 ( .B1(n8757), .B2(n9368), .C1(n8733), .C2(n9365), .A(n1815), 
        .ZN(n1812) );
  AOI22_X1 U1738 ( .A1(n9362), .A2(n10090), .B1(n9359), .B2(n10122), .ZN(n1815) );
  OAI221_X1 U1739 ( .B1(n8391), .B2(n9428), .C1(n8359), .C2(n9425), .A(n1788), 
        .ZN(n1787) );
  AOI22_X1 U1740 ( .A1(n9422), .A2(n10641), .B1(n9419), .B2(n10521), .ZN(n1788) );
  OAI221_X1 U1741 ( .B1(n8758), .B2(n9368), .C1(n8734), .C2(n9365), .A(n1797), 
        .ZN(n1794) );
  AOI22_X1 U1742 ( .A1(n9362), .A2(n10089), .B1(n9359), .B2(n10121), .ZN(n1797) );
  OAI221_X1 U1743 ( .B1(n8392), .B2(n9428), .C1(n8360), .C2(n9425), .A(n1770), 
        .ZN(n1769) );
  AOI22_X1 U1744 ( .A1(n9422), .A2(n10640), .B1(n9419), .B2(n10520), .ZN(n1770) );
  OAI221_X1 U1745 ( .B1(n8759), .B2(n9368), .C1(n8735), .C2(n9365), .A(n1779), 
        .ZN(n1776) );
  AOI22_X1 U1746 ( .A1(n9362), .A2(n10088), .B1(n9359), .B2(n10120), .ZN(n1779) );
  OAI221_X1 U1747 ( .B1(n8393), .B2(n9428), .C1(n8361), .C2(n9425), .A(n1752), 
        .ZN(n1751) );
  AOI22_X1 U1748 ( .A1(n9422), .A2(n10639), .B1(n9419), .B2(n10519), .ZN(n1752) );
  OAI221_X1 U1749 ( .B1(n8760), .B2(n9368), .C1(n8736), .C2(n9365), .A(n1761), 
        .ZN(n1758) );
  AOI22_X1 U1750 ( .A1(n9362), .A2(n10087), .B1(n9359), .B2(n10119), .ZN(n1761) );
  OAI221_X1 U1751 ( .B1(n8394), .B2(n9428), .C1(n8362), .C2(n9425), .A(n1734), 
        .ZN(n1733) );
  AOI22_X1 U1752 ( .A1(n9422), .A2(n10638), .B1(n9419), .B2(n10518), .ZN(n1734) );
  OAI221_X1 U1753 ( .B1(n8761), .B2(n9368), .C1(n8737), .C2(n9365), .A(n1743), 
        .ZN(n1740) );
  AOI22_X1 U1754 ( .A1(n9362), .A2(n10086), .B1(n9359), .B2(n10118), .ZN(n1743) );
  OAI221_X1 U1755 ( .B1(n8395), .B2(n9428), .C1(n8363), .C2(n9425), .A(n1716), 
        .ZN(n1715) );
  AOI22_X1 U1756 ( .A1(n9422), .A2(n10637), .B1(n9418), .B2(n10517), .ZN(n1716) );
  OAI221_X1 U1757 ( .B1(n8762), .B2(n9368), .C1(n8738), .C2(n9365), .A(n1725), 
        .ZN(n1722) );
  AOI22_X1 U1758 ( .A1(n9362), .A2(n10085), .B1(n9358), .B2(n10117), .ZN(n1725) );
  OAI221_X1 U1759 ( .B1(n8396), .B2(n9428), .C1(n8364), .C2(n9425), .A(n1698), 
        .ZN(n1697) );
  AOI22_X1 U1760 ( .A1(n9422), .A2(n10636), .B1(n9418), .B2(n10516), .ZN(n1698) );
  OAI221_X1 U1761 ( .B1(n8763), .B2(n9368), .C1(n8739), .C2(n9365), .A(n1707), 
        .ZN(n1704) );
  AOI22_X1 U1762 ( .A1(n9362), .A2(n10084), .B1(n9358), .B2(n10116), .ZN(n1707) );
  OAI221_X1 U1763 ( .B1(n8397), .B2(n9428), .C1(n8365), .C2(n9425), .A(n1680), 
        .ZN(n1679) );
  AOI22_X1 U1764 ( .A1(n9422), .A2(n10635), .B1(n9418), .B2(n10515), .ZN(n1680) );
  OAI221_X1 U1765 ( .B1(n8764), .B2(n9368), .C1(n8740), .C2(n9365), .A(n1689), 
        .ZN(n1686) );
  AOI22_X1 U1766 ( .A1(n9362), .A2(n10083), .B1(n9358), .B2(n10115), .ZN(n1689) );
  OAI221_X1 U1767 ( .B1(n8398), .B2(n9428), .C1(n8366), .C2(n9425), .A(n1662), 
        .ZN(n1661) );
  AOI22_X1 U1768 ( .A1(n9422), .A2(n10634), .B1(n9418), .B2(n10514), .ZN(n1662) );
  OAI221_X1 U1769 ( .B1(n8765), .B2(n9368), .C1(n8741), .C2(n9365), .A(n1671), 
        .ZN(n1668) );
  AOI22_X1 U1770 ( .A1(n9362), .A2(n10082), .B1(n9358), .B2(n10114), .ZN(n1671) );
  OAI221_X1 U1771 ( .B1(n8399), .B2(n9429), .C1(n8367), .C2(n9426), .A(n1644), 
        .ZN(n1643) );
  AOI22_X1 U1772 ( .A1(n9423), .A2(n10561), .B1(n9418), .B2(n10513), .ZN(n1644) );
  OAI221_X1 U1773 ( .B1(n8766), .B2(n9369), .C1(n8287), .C2(n9366), .A(n1653), 
        .ZN(n1650) );
  AOI22_X1 U1774 ( .A1(n9363), .A2(n10081), .B1(n9358), .B2(n10113), .ZN(n1653) );
  OAI221_X1 U1775 ( .B1(n8400), .B2(n9429), .C1(n8368), .C2(n9426), .A(n1626), 
        .ZN(n1625) );
  AOI22_X1 U1776 ( .A1(n9423), .A2(n10560), .B1(n9418), .B2(n10512), .ZN(n1626) );
  OAI221_X1 U1777 ( .B1(n8767), .B2(n9369), .C1(n8288), .C2(n9366), .A(n1635), 
        .ZN(n1632) );
  AOI22_X1 U1778 ( .A1(n9363), .A2(n10080), .B1(n9358), .B2(n10112), .ZN(n1635) );
  OAI221_X1 U1779 ( .B1(n8401), .B2(n9429), .C1(n8369), .C2(n9426), .A(n1608), 
        .ZN(n1607) );
  AOI22_X1 U1780 ( .A1(n9423), .A2(n10559), .B1(n9418), .B2(n10511), .ZN(n1608) );
  OAI221_X1 U1781 ( .B1(n8768), .B2(n9369), .C1(n8289), .C2(n9366), .A(n1617), 
        .ZN(n1614) );
  AOI22_X1 U1782 ( .A1(n9363), .A2(n10079), .B1(n9358), .B2(n10111), .ZN(n1617) );
  OAI221_X1 U1783 ( .B1(n8402), .B2(n9429), .C1(n8370), .C2(n9426), .A(n1590), 
        .ZN(n1589) );
  AOI22_X1 U1784 ( .A1(n9423), .A2(n10558), .B1(n9418), .B2(n10510), .ZN(n1590) );
  OAI221_X1 U1785 ( .B1(n8769), .B2(n9369), .C1(n8290), .C2(n9366), .A(n1599), 
        .ZN(n1596) );
  AOI22_X1 U1786 ( .A1(n9363), .A2(n10078), .B1(n9358), .B2(n10110), .ZN(n1599) );
  OAI221_X1 U1787 ( .B1(n8403), .B2(n9429), .C1(n8371), .C2(n9426), .A(n1572), 
        .ZN(n1571) );
  AOI22_X1 U1788 ( .A1(n9423), .A2(n10557), .B1(n9418), .B2(n10509), .ZN(n1572) );
  OAI221_X1 U1789 ( .B1(n8770), .B2(n9369), .C1(n8291), .C2(n9366), .A(n1581), 
        .ZN(n1578) );
  AOI22_X1 U1790 ( .A1(n9363), .A2(n10077), .B1(n9358), .B2(n10109), .ZN(n1581) );
  OAI221_X1 U1791 ( .B1(n8404), .B2(n9429), .C1(n8372), .C2(n9426), .A(n1554), 
        .ZN(n1553) );
  AOI22_X1 U1792 ( .A1(n9423), .A2(n10556), .B1(n9418), .B2(n10508), .ZN(n1554) );
  OAI221_X1 U1793 ( .B1(n8771), .B2(n9369), .C1(n8292), .C2(n9366), .A(n1563), 
        .ZN(n1560) );
  AOI22_X1 U1794 ( .A1(n9363), .A2(n10076), .B1(n9358), .B2(n10108), .ZN(n1563) );
  OAI221_X1 U1795 ( .B1(n8405), .B2(n9429), .C1(n8373), .C2(n9426), .A(n1536), 
        .ZN(n1535) );
  AOI22_X1 U1796 ( .A1(n9423), .A2(n10555), .B1(n9418), .B2(n10507), .ZN(n1536) );
  OAI221_X1 U1797 ( .B1(n8772), .B2(n9369), .C1(n8293), .C2(n9366), .A(n1545), 
        .ZN(n1542) );
  AOI22_X1 U1798 ( .A1(n9363), .A2(n10075), .B1(n9358), .B2(n10107), .ZN(n1545) );
  OAI221_X1 U1799 ( .B1(n8406), .B2(n9429), .C1(n8374), .C2(n9426), .A(n1488), 
        .ZN(n1485) );
  AOI22_X1 U1800 ( .A1(n9423), .A2(n10554), .B1(n9418), .B2(n10506), .ZN(n1488) );
  OAI221_X1 U1801 ( .B1(n8773), .B2(n9369), .C1(n8294), .C2(n9366), .A(n1517), 
        .ZN(n1508) );
  AOI22_X1 U1802 ( .A1(n9363), .A2(n10074), .B1(n9358), .B2(n10106), .ZN(n1517) );
  OAI22_X1 U1803 ( .A1(n9329), .A2(n9603), .B1(n8655), .B2(n9612), .ZN(n3199)
         );
  OAI22_X1 U1804 ( .A1(n9326), .A2(n9603), .B1(n8656), .B2(n9612), .ZN(n3200)
         );
  OAI22_X1 U1805 ( .A1(n9323), .A2(n9603), .B1(n8657), .B2(n9612), .ZN(n3201)
         );
  OAI22_X1 U1806 ( .A1(n9320), .A2(n9603), .B1(n8658), .B2(n9611), .ZN(n3202)
         );
  OAI22_X1 U1807 ( .A1(n9317), .A2(n9603), .B1(n8659), .B2(n9611), .ZN(n3203)
         );
  OAI22_X1 U1808 ( .A1(n9311), .A2(n9603), .B1(n8661), .B2(n9611), .ZN(n3205)
         );
  OAI22_X1 U1809 ( .A1(n9308), .A2(n9603), .B1(n8662), .B2(n9610), .ZN(n3206)
         );
  OAI22_X1 U1810 ( .A1(n9305), .A2(n9603), .B1(n8663), .B2(n9610), .ZN(n3207)
         );
  OAI22_X1 U1811 ( .A1(n9302), .A2(n9603), .B1(n8664), .B2(n9610), .ZN(n3208)
         );
  OAI22_X1 U1812 ( .A1(n9299), .A2(n9603), .B1(n8665), .B2(n9610), .ZN(n3209)
         );
  OAI22_X1 U1813 ( .A1(n9296), .A2(n9604), .B1(n8666), .B2(n9609), .ZN(n3210)
         );
  OAI22_X1 U1814 ( .A1(n9290), .A2(n9604), .B1(n8668), .B2(n9609), .ZN(n3212)
         );
  OAI22_X1 U1815 ( .A1(n9287), .A2(n9604), .B1(n8669), .B2(n9609), .ZN(n3213)
         );
  OAI22_X1 U1816 ( .A1(n9284), .A2(n9604), .B1(n8670), .B2(n9608), .ZN(n3214)
         );
  OAI22_X1 U1817 ( .A1(n9278), .A2(n9604), .B1(n8672), .B2(n9608), .ZN(n3216)
         );
  OAI22_X1 U1818 ( .A1(n9275), .A2(n9604), .B1(n8673), .B2(n9608), .ZN(n3217)
         );
  OAI22_X1 U1819 ( .A1(n9272), .A2(n9604), .B1(n8674), .B2(n9607), .ZN(n3218)
         );
  OAI22_X1 U1820 ( .A1(n9269), .A2(n9604), .B1(n8675), .B2(n9607), .ZN(n3219)
         );
  OAI22_X1 U1821 ( .A1(n9266), .A2(n9604), .B1(n8676), .B2(n9607), .ZN(n3220)
         );
  OAI22_X1 U1822 ( .A1(n9263), .A2(n9604), .B1(n8677), .B2(n9607), .ZN(n3221)
         );
  OAI22_X1 U1823 ( .A1(n9260), .A2(n9603), .B1(n8678), .B2(n9606), .ZN(n3222)
         );
  OAI22_X1 U1824 ( .A1(n9257), .A2(n9604), .B1(n8679), .B2(n9606), .ZN(n3223)
         );
  OAI22_X1 U1825 ( .A1(n9254), .A2(n9603), .B1(n8680), .B2(n9606), .ZN(n3224)
         );
  OAI22_X1 U1826 ( .A1(n9251), .A2(n9604), .B1(n8681), .B2(n9606), .ZN(n3225)
         );
  OAI22_X1 U1827 ( .A1(n9248), .A2(n9603), .B1(n8682), .B2(n9605), .ZN(n3226)
         );
  OAI22_X1 U1828 ( .A1(n9245), .A2(n9604), .B1(n8683), .B2(n9605), .ZN(n3227)
         );
  OAI22_X1 U1829 ( .A1(n9242), .A2(n9603), .B1(n8684), .B2(n9605), .ZN(n3228)
         );
  OAI22_X1 U1830 ( .A1(n9239), .A2(n9604), .B1(n8685), .B2(n9605), .ZN(n3229)
         );
  OAI22_X1 U1831 ( .A1(n9331), .A2(n9835), .B1(n2351), .B2(n9836), .ZN(n9109)
         );
  OAI22_X1 U1832 ( .A1(n9328), .A2(n9834), .B1(n2343), .B2(n9836), .ZN(n9108)
         );
  OAI22_X1 U1833 ( .A1(n9325), .A2(n9835), .B1(n2335), .B2(n9836), .ZN(n9107)
         );
  OAI22_X1 U1834 ( .A1(n9322), .A2(n9834), .B1(n2327), .B2(n9836), .ZN(n9106)
         );
  OAI22_X1 U1835 ( .A1(n9319), .A2(n9835), .B1(n2319), .B2(n9837), .ZN(n9105)
         );
  OAI22_X1 U1836 ( .A1(n9316), .A2(n9834), .B1(n2311), .B2(n9837), .ZN(n9104)
         );
  OAI22_X1 U1837 ( .A1(n9313), .A2(n9835), .B1(n2303), .B2(n9837), .ZN(n9103)
         );
  OAI22_X1 U1838 ( .A1(n9310), .A2(n9834), .B1(n2295), .B2(n9837), .ZN(n9102)
         );
  OAI22_X1 U1839 ( .A1(n9307), .A2(n9835), .B1(n2287), .B2(n9838), .ZN(n9101)
         );
  OAI22_X1 U1840 ( .A1(n9304), .A2(n9835), .B1(n2279), .B2(n9838), .ZN(n9100)
         );
  OAI22_X1 U1841 ( .A1(n9301), .A2(n9835), .B1(n2271), .B2(n9838), .ZN(n9099)
         );
  OAI22_X1 U1842 ( .A1(n9298), .A2(n9835), .B1(n2263), .B2(n9838), .ZN(n9098)
         );
  OAI22_X1 U1843 ( .A1(n9295), .A2(n9835), .B1(n2255), .B2(n9839), .ZN(n9097)
         );
  OAI22_X1 U1844 ( .A1(n9292), .A2(n9835), .B1(n2247), .B2(n9839), .ZN(n9096)
         );
  OAI22_X1 U1845 ( .A1(n9289), .A2(n9835), .B1(n2239), .B2(n9839), .ZN(n9095)
         );
  OAI22_X1 U1846 ( .A1(n9286), .A2(n9835), .B1(n2231), .B2(n9839), .ZN(n9094)
         );
  OAI22_X1 U1847 ( .A1(n9283), .A2(n9835), .B1(n2223), .B2(n9840), .ZN(n9093)
         );
  OAI22_X1 U1848 ( .A1(n9280), .A2(n9835), .B1(n2215), .B2(n9840), .ZN(n9092)
         );
  OAI22_X1 U1849 ( .A1(n9277), .A2(n9835), .B1(n2207), .B2(n9840), .ZN(n9091)
         );
  OAI22_X1 U1850 ( .A1(n9274), .A2(n9835), .B1(n2199), .B2(n9840), .ZN(n9090)
         );
  OAI22_X1 U1851 ( .A1(n9271), .A2(n9834), .B1(n2191), .B2(n9841), .ZN(n9089)
         );
  OAI22_X1 U1852 ( .A1(n9268), .A2(n9834), .B1(n2183), .B2(n9841), .ZN(n9088)
         );
  OAI22_X1 U1853 ( .A1(n9265), .A2(n9834), .B1(n2175), .B2(n9841), .ZN(n9087)
         );
  OAI22_X1 U1854 ( .A1(n9262), .A2(n9834), .B1(n2167), .B2(n9841), .ZN(n9086)
         );
  OAI22_X1 U1855 ( .A1(n9259), .A2(n9834), .B1(n2159), .B2(n9842), .ZN(n9085)
         );
  OAI22_X1 U1856 ( .A1(n9256), .A2(n9834), .B1(n2151), .B2(n9842), .ZN(n9084)
         );
  OAI22_X1 U1857 ( .A1(n9253), .A2(n9834), .B1(n2143), .B2(n9842), .ZN(n9083)
         );
  OAI22_X1 U1858 ( .A1(n9250), .A2(n9834), .B1(n2135), .B2(n9842), .ZN(n9082)
         );
  OAI22_X1 U1859 ( .A1(n9247), .A2(n9834), .B1(n2127), .B2(n9843), .ZN(n9081)
         );
  OAI22_X1 U1860 ( .A1(n9244), .A2(n9834), .B1(n2119), .B2(n9843), .ZN(n9080)
         );
  OAI22_X1 U1861 ( .A1(n9241), .A2(n9834), .B1(n2111), .B2(n9843), .ZN(n9079)
         );
  OAI22_X1 U1862 ( .A1(n9238), .A2(n9834), .B1(n2103), .B2(n9843), .ZN(n9078)
         );
  OAI22_X1 U1863 ( .A1(n9331), .A2(n9747), .B1(n8439), .B2(n9748), .ZN(n3955)
         );
  OAI22_X1 U1864 ( .A1(n9328), .A2(n9746), .B1(n8440), .B2(n9748), .ZN(n3939)
         );
  OAI22_X1 U1865 ( .A1(n9325), .A2(n9747), .B1(n8441), .B2(n9748), .ZN(n3923)
         );
  OAI22_X1 U1866 ( .A1(n9322), .A2(n9746), .B1(n8442), .B2(n9748), .ZN(n3907)
         );
  OAI22_X1 U1867 ( .A1(n9319), .A2(n9747), .B1(n8443), .B2(n9749), .ZN(n3891)
         );
  OAI22_X1 U1868 ( .A1(n9316), .A2(n9746), .B1(n8444), .B2(n9749), .ZN(n3875)
         );
  OAI22_X1 U1869 ( .A1(n9313), .A2(n9747), .B1(n8445), .B2(n9749), .ZN(n3859)
         );
  OAI22_X1 U1870 ( .A1(n9310), .A2(n9746), .B1(n8446), .B2(n9749), .ZN(n3843)
         );
  OAI22_X1 U1871 ( .A1(n9307), .A2(n9747), .B1(n8447), .B2(n9750), .ZN(n3827)
         );
  OAI22_X1 U1872 ( .A1(n9304), .A2(n9747), .B1(n8448), .B2(n9750), .ZN(n3811)
         );
  OAI22_X1 U1873 ( .A1(n9301), .A2(n9747), .B1(n8449), .B2(n9750), .ZN(n3795)
         );
  OAI22_X1 U1874 ( .A1(n9298), .A2(n9747), .B1(n8450), .B2(n9750), .ZN(n3779)
         );
  OAI22_X1 U1875 ( .A1(n9295), .A2(n9747), .B1(n8451), .B2(n9751), .ZN(n3763)
         );
  OAI22_X1 U1876 ( .A1(n9292), .A2(n9747), .B1(n8452), .B2(n9751), .ZN(n3747)
         );
  OAI22_X1 U1877 ( .A1(n9289), .A2(n9747), .B1(n8453), .B2(n9751), .ZN(n3731)
         );
  OAI22_X1 U1878 ( .A1(n9286), .A2(n9747), .B1(n8454), .B2(n9751), .ZN(n3715)
         );
  OAI22_X1 U1879 ( .A1(n9283), .A2(n9747), .B1(n8455), .B2(n9752), .ZN(n3699)
         );
  OAI22_X1 U1880 ( .A1(n9280), .A2(n9747), .B1(n8456), .B2(n9752), .ZN(n3683)
         );
  OAI22_X1 U1881 ( .A1(n9277), .A2(n9747), .B1(n8457), .B2(n9752), .ZN(n3667)
         );
  OAI22_X1 U1882 ( .A1(n9274), .A2(n9747), .B1(n8458), .B2(n9752), .ZN(n3651)
         );
  OAI22_X1 U1883 ( .A1(n9271), .A2(n9746), .B1(n8459), .B2(n9753), .ZN(n3635)
         );
  OAI22_X1 U1884 ( .A1(n9268), .A2(n9746), .B1(n8460), .B2(n9753), .ZN(n3619)
         );
  OAI22_X1 U1885 ( .A1(n9265), .A2(n9746), .B1(n8461), .B2(n9753), .ZN(n3603)
         );
  OAI22_X1 U1886 ( .A1(n9262), .A2(n9746), .B1(n8462), .B2(n9753), .ZN(n3587)
         );
  OAI22_X1 U1887 ( .A1(n9259), .A2(n9746), .B1(n8463), .B2(n9754), .ZN(n3571)
         );
  OAI22_X1 U1888 ( .A1(n9256), .A2(n9746), .B1(n8464), .B2(n9754), .ZN(n3555)
         );
  OAI22_X1 U1889 ( .A1(n9253), .A2(n9746), .B1(n8465), .B2(n9754), .ZN(n3539)
         );
  OAI22_X1 U1890 ( .A1(n9250), .A2(n9746), .B1(n8466), .B2(n9754), .ZN(n3523)
         );
  OAI22_X1 U1891 ( .A1(n9247), .A2(n9746), .B1(n8467), .B2(n9755), .ZN(n3507)
         );
  OAI22_X1 U1892 ( .A1(n9244), .A2(n9746), .B1(n8468), .B2(n9755), .ZN(n3491)
         );
  OAI22_X1 U1893 ( .A1(n9241), .A2(n9746), .B1(n8469), .B2(n9755), .ZN(n3475)
         );
  OAI22_X1 U1894 ( .A1(n9238), .A2(n9746), .B1(n8470), .B2(n9755), .ZN(n3459)
         );
  OAI22_X1 U1895 ( .A1(n9331), .A2(n9736), .B1(n8510), .B2(n9737), .ZN(n3954)
         );
  OAI22_X1 U1896 ( .A1(n9328), .A2(n9735), .B1(n8511), .B2(n9737), .ZN(n3938)
         );
  OAI22_X1 U1897 ( .A1(n9325), .A2(n9736), .B1(n8512), .B2(n9737), .ZN(n3922)
         );
  OAI22_X1 U1898 ( .A1(n9322), .A2(n9735), .B1(n8513), .B2(n9737), .ZN(n3906)
         );
  OAI22_X1 U1899 ( .A1(n9319), .A2(n9736), .B1(n8514), .B2(n9738), .ZN(n3890)
         );
  OAI22_X1 U1900 ( .A1(n9316), .A2(n9735), .B1(n8515), .B2(n9738), .ZN(n3874)
         );
  OAI22_X1 U1901 ( .A1(n9313), .A2(n9736), .B1(n8516), .B2(n9738), .ZN(n3858)
         );
  OAI22_X1 U1902 ( .A1(n9310), .A2(n9735), .B1(n8517), .B2(n9738), .ZN(n3842)
         );
  OAI22_X1 U1903 ( .A1(n9307), .A2(n9736), .B1(n8518), .B2(n9739), .ZN(n3826)
         );
  OAI22_X1 U1904 ( .A1(n9304), .A2(n9736), .B1(n8519), .B2(n9739), .ZN(n3810)
         );
  OAI22_X1 U1905 ( .A1(n9301), .A2(n9736), .B1(n8520), .B2(n9739), .ZN(n3794)
         );
  OAI22_X1 U1906 ( .A1(n9298), .A2(n9736), .B1(n8521), .B2(n9739), .ZN(n3778)
         );
  OAI22_X1 U1907 ( .A1(n9295), .A2(n9736), .B1(n8522), .B2(n9740), .ZN(n3762)
         );
  OAI22_X1 U1908 ( .A1(n9292), .A2(n9736), .B1(n8523), .B2(n9740), .ZN(n3746)
         );
  OAI22_X1 U1909 ( .A1(n9289), .A2(n9736), .B1(n8524), .B2(n9740), .ZN(n3730)
         );
  OAI22_X1 U1910 ( .A1(n9286), .A2(n9736), .B1(n8525), .B2(n9740), .ZN(n3714)
         );
  OAI22_X1 U1911 ( .A1(n9283), .A2(n9736), .B1(n8526), .B2(n9741), .ZN(n3698)
         );
  OAI22_X1 U1912 ( .A1(n9280), .A2(n9736), .B1(n8527), .B2(n9741), .ZN(n3682)
         );
  OAI22_X1 U1913 ( .A1(n9277), .A2(n9736), .B1(n8528), .B2(n9741), .ZN(n3666)
         );
  OAI22_X1 U1914 ( .A1(n9274), .A2(n9736), .B1(n8529), .B2(n9741), .ZN(n3650)
         );
  OAI22_X1 U1915 ( .A1(n9271), .A2(n9735), .B1(n8530), .B2(n9742), .ZN(n3634)
         );
  OAI22_X1 U1916 ( .A1(n9268), .A2(n9735), .B1(n8531), .B2(n9742), .ZN(n3618)
         );
  OAI22_X1 U1917 ( .A1(n9265), .A2(n9735), .B1(n8532), .B2(n9742), .ZN(n3602)
         );
  OAI22_X1 U1918 ( .A1(n9262), .A2(n9735), .B1(n8533), .B2(n9742), .ZN(n3586)
         );
  OAI22_X1 U1919 ( .A1(n9259), .A2(n9735), .B1(n8534), .B2(n9743), .ZN(n3570)
         );
  OAI22_X1 U1920 ( .A1(n9256), .A2(n9735), .B1(n8535), .B2(n9743), .ZN(n3554)
         );
  OAI22_X1 U1921 ( .A1(n9253), .A2(n9735), .B1(n8536), .B2(n9743), .ZN(n3538)
         );
  OAI22_X1 U1922 ( .A1(n9250), .A2(n9735), .B1(n8537), .B2(n9743), .ZN(n3522)
         );
  OAI22_X1 U1923 ( .A1(n9247), .A2(n9735), .B1(n8538), .B2(n9744), .ZN(n3506)
         );
  OAI22_X1 U1924 ( .A1(n9244), .A2(n9735), .B1(n8539), .B2(n9744), .ZN(n3490)
         );
  OAI22_X1 U1925 ( .A1(n9241), .A2(n9735), .B1(n8540), .B2(n9744), .ZN(n3474)
         );
  OAI22_X1 U1926 ( .A1(n9238), .A2(n9735), .B1(n8541), .B2(n9744), .ZN(n3458)
         );
  OAI22_X1 U1927 ( .A1(n9329), .A2(n9725), .B1(n8599), .B2(n9726), .ZN(n3936)
         );
  OAI22_X1 U1928 ( .A1(n9326), .A2(n9724), .B1(n8600), .B2(n9726), .ZN(n3920)
         );
  OAI22_X1 U1929 ( .A1(n9323), .A2(n9725), .B1(n8601), .B2(n9726), .ZN(n3904)
         );
  OAI22_X1 U1930 ( .A1(n9320), .A2(n9724), .B1(n8602), .B2(n9727), .ZN(n3888)
         );
  OAI22_X1 U1931 ( .A1(n9317), .A2(n9725), .B1(n8603), .B2(n9727), .ZN(n3872)
         );
  OAI22_X1 U1932 ( .A1(n9314), .A2(n9724), .B1(n8604), .B2(n9727), .ZN(n3856)
         );
  OAI22_X1 U1933 ( .A1(n9311), .A2(n9725), .B1(n8605), .B2(n9727), .ZN(n3840)
         );
  OAI22_X1 U1934 ( .A1(n9308), .A2(n9725), .B1(n8606), .B2(n9728), .ZN(n3824)
         );
  OAI22_X1 U1935 ( .A1(n9305), .A2(n9725), .B1(n8607), .B2(n9728), .ZN(n3808)
         );
  OAI22_X1 U1936 ( .A1(n9302), .A2(n9725), .B1(n8608), .B2(n9728), .ZN(n3792)
         );
  OAI22_X1 U1937 ( .A1(n9299), .A2(n9725), .B1(n8609), .B2(n9728), .ZN(n3776)
         );
  OAI22_X1 U1938 ( .A1(n9296), .A2(n9725), .B1(n8610), .B2(n9729), .ZN(n3760)
         );
  OAI22_X1 U1939 ( .A1(n9293), .A2(n9725), .B1(n8611), .B2(n9729), .ZN(n3744)
         );
  OAI22_X1 U1940 ( .A1(n9290), .A2(n9725), .B1(n8612), .B2(n9729), .ZN(n3728)
         );
  OAI22_X1 U1941 ( .A1(n9287), .A2(n9725), .B1(n8613), .B2(n9729), .ZN(n3712)
         );
  OAI22_X1 U1942 ( .A1(n9284), .A2(n9725), .B1(n8614), .B2(n9730), .ZN(n3696)
         );
  OAI22_X1 U1943 ( .A1(n9281), .A2(n9725), .B1(n8615), .B2(n9730), .ZN(n3680)
         );
  OAI22_X1 U1944 ( .A1(n9278), .A2(n9725), .B1(n8616), .B2(n9730), .ZN(n3664)
         );
  OAI22_X1 U1945 ( .A1(n9275), .A2(n9725), .B1(n8617), .B2(n9730), .ZN(n3648)
         );
  OAI22_X1 U1946 ( .A1(n9272), .A2(n9724), .B1(n8618), .B2(n9731), .ZN(n3632)
         );
  OAI22_X1 U1947 ( .A1(n9269), .A2(n9724), .B1(n8619), .B2(n9731), .ZN(n3616)
         );
  OAI22_X1 U1948 ( .A1(n9266), .A2(n9724), .B1(n8620), .B2(n9731), .ZN(n3600)
         );
  OAI22_X1 U1949 ( .A1(n9263), .A2(n9724), .B1(n8621), .B2(n9731), .ZN(n3584)
         );
  OAI22_X1 U1950 ( .A1(n9260), .A2(n9724), .B1(n8622), .B2(n9732), .ZN(n3568)
         );
  OAI22_X1 U1951 ( .A1(n9257), .A2(n9724), .B1(n8623), .B2(n9732), .ZN(n3552)
         );
  OAI22_X1 U1952 ( .A1(n9254), .A2(n9724), .B1(n8624), .B2(n9732), .ZN(n3536)
         );
  OAI22_X1 U1953 ( .A1(n9251), .A2(n9724), .B1(n8625), .B2(n9732), .ZN(n3520)
         );
  OAI22_X1 U1954 ( .A1(n9248), .A2(n9724), .B1(n8626), .B2(n9733), .ZN(n3504)
         );
  OAI22_X1 U1955 ( .A1(n9245), .A2(n9724), .B1(n8627), .B2(n9733), .ZN(n3488)
         );
  OAI22_X1 U1956 ( .A1(n9242), .A2(n9724), .B1(n8628), .B2(n9733), .ZN(n3472)
         );
  OAI22_X1 U1957 ( .A1(n9239), .A2(n9724), .B1(n8629), .B2(n9733), .ZN(n3456)
         );
  OAI22_X1 U1958 ( .A1(n9332), .A2(n9625), .B1(n8742), .B2(n9634), .ZN(n3262)
         );
  OAI22_X1 U1959 ( .A1(n9329), .A2(n9625), .B1(n8743), .B2(n9634), .ZN(n3263)
         );
  OAI22_X1 U1960 ( .A1(n9326), .A2(n9625), .B1(n8744), .B2(n9634), .ZN(n3264)
         );
  OAI22_X1 U1961 ( .A1(n9323), .A2(n9625), .B1(n8745), .B2(n9634), .ZN(n3265)
         );
  OAI22_X1 U1962 ( .A1(n9320), .A2(n9625), .B1(n8746), .B2(n9633), .ZN(n3266)
         );
  OAI22_X1 U1963 ( .A1(n9317), .A2(n9625), .B1(n8747), .B2(n9633), .ZN(n3267)
         );
  OAI22_X1 U1964 ( .A1(n9314), .A2(n9625), .B1(n8748), .B2(n9633), .ZN(n3268)
         );
  OAI22_X1 U1965 ( .A1(n9311), .A2(n9625), .B1(n8749), .B2(n9633), .ZN(n3269)
         );
  OAI22_X1 U1966 ( .A1(n9308), .A2(n9625), .B1(n8750), .B2(n9632), .ZN(n3270)
         );
  OAI22_X1 U1967 ( .A1(n9305), .A2(n9625), .B1(n8751), .B2(n9632), .ZN(n3271)
         );
  OAI22_X1 U1968 ( .A1(n9302), .A2(n9625), .B1(n8752), .B2(n9632), .ZN(n3272)
         );
  OAI22_X1 U1969 ( .A1(n9299), .A2(n9625), .B1(n8753), .B2(n9632), .ZN(n3273)
         );
  OAI22_X1 U1970 ( .A1(n9296), .A2(n9626), .B1(n8754), .B2(n9631), .ZN(n3274)
         );
  OAI22_X1 U1971 ( .A1(n9293), .A2(n9626), .B1(n8755), .B2(n9631), .ZN(n3275)
         );
  OAI22_X1 U1972 ( .A1(n9290), .A2(n9626), .B1(n8756), .B2(n9631), .ZN(n3276)
         );
  OAI22_X1 U1973 ( .A1(n9287), .A2(n9626), .B1(n8757), .B2(n9631), .ZN(n3277)
         );
  OAI22_X1 U1974 ( .A1(n9284), .A2(n9626), .B1(n8758), .B2(n9630), .ZN(n3278)
         );
  OAI22_X1 U1975 ( .A1(n9281), .A2(n9626), .B1(n8759), .B2(n9630), .ZN(n3279)
         );
  OAI22_X1 U1976 ( .A1(n9278), .A2(n9626), .B1(n8760), .B2(n9630), .ZN(n3280)
         );
  OAI22_X1 U1977 ( .A1(n9275), .A2(n9626), .B1(n8761), .B2(n9630), .ZN(n3281)
         );
  OAI22_X1 U1978 ( .A1(n9272), .A2(n9626), .B1(n8762), .B2(n9629), .ZN(n3282)
         );
  OAI22_X1 U1979 ( .A1(n9269), .A2(n9626), .B1(n8763), .B2(n9629), .ZN(n3283)
         );
  OAI22_X1 U1980 ( .A1(n9266), .A2(n9626), .B1(n8764), .B2(n9629), .ZN(n3284)
         );
  OAI22_X1 U1981 ( .A1(n9263), .A2(n9626), .B1(n8765), .B2(n9629), .ZN(n3285)
         );
  OAI22_X1 U1982 ( .A1(n9260), .A2(n9625), .B1(n8766), .B2(n9628), .ZN(n3286)
         );
  OAI22_X1 U1983 ( .A1(n9257), .A2(n9626), .B1(n8767), .B2(n9628), .ZN(n3287)
         );
  OAI22_X1 U1984 ( .A1(n9254), .A2(n9625), .B1(n8768), .B2(n9628), .ZN(n3288)
         );
  OAI22_X1 U1985 ( .A1(n9251), .A2(n9626), .B1(n8769), .B2(n9628), .ZN(n3289)
         );
  OAI22_X1 U1986 ( .A1(n9248), .A2(n9625), .B1(n8770), .B2(n9627), .ZN(n3290)
         );
  OAI22_X1 U1987 ( .A1(n9245), .A2(n9626), .B1(n8771), .B2(n9627), .ZN(n3291)
         );
  OAI22_X1 U1988 ( .A1(n9242), .A2(n9625), .B1(n8772), .B2(n9627), .ZN(n3292)
         );
  OAI22_X1 U1989 ( .A1(n9239), .A2(n9626), .B1(n8773), .B2(n9627), .ZN(n3293)
         );
  OAI22_X1 U1990 ( .A1(n9332), .A2(n9692), .B1(n8830), .B2(n9693), .ZN(n3946)
         );
  OAI22_X1 U1991 ( .A1(n9329), .A2(n9691), .B1(n8831), .B2(n9693), .ZN(n3930)
         );
  OAI22_X1 U1992 ( .A1(n9326), .A2(n9692), .B1(n8832), .B2(n9693), .ZN(n3914)
         );
  OAI22_X1 U1993 ( .A1(n9323), .A2(n9691), .B1(n8833), .B2(n9693), .ZN(n3898)
         );
  OAI22_X1 U1994 ( .A1(n9320), .A2(n9692), .B1(n8834), .B2(n9694), .ZN(n3882)
         );
  OAI22_X1 U1995 ( .A1(n9317), .A2(n9691), .B1(n8835), .B2(n9694), .ZN(n3866)
         );
  OAI22_X1 U1996 ( .A1(n9314), .A2(n9692), .B1(n8836), .B2(n9694), .ZN(n3850)
         );
  OAI22_X1 U1997 ( .A1(n9311), .A2(n9691), .B1(n8837), .B2(n9694), .ZN(n3834)
         );
  OAI22_X1 U1998 ( .A1(n9308), .A2(n9692), .B1(n8838), .B2(n9695), .ZN(n3818)
         );
  OAI22_X1 U1999 ( .A1(n9305), .A2(n9692), .B1(n8839), .B2(n9695), .ZN(n3802)
         );
  OAI22_X1 U2000 ( .A1(n9302), .A2(n9692), .B1(n8840), .B2(n9695), .ZN(n3786)
         );
  OAI22_X1 U2001 ( .A1(n9299), .A2(n9692), .B1(n8841), .B2(n9695), .ZN(n3770)
         );
  OAI22_X1 U2002 ( .A1(n9296), .A2(n9692), .B1(n8842), .B2(n9696), .ZN(n3754)
         );
  OAI22_X1 U2003 ( .A1(n9293), .A2(n9692), .B1(n8843), .B2(n9696), .ZN(n3738)
         );
  OAI22_X1 U2004 ( .A1(n9290), .A2(n9692), .B1(n8844), .B2(n9696), .ZN(n3722)
         );
  OAI22_X1 U2005 ( .A1(n9287), .A2(n9692), .B1(n8845), .B2(n9696), .ZN(n3706)
         );
  OAI22_X1 U2006 ( .A1(n9284), .A2(n9692), .B1(n8846), .B2(n9697), .ZN(n3690)
         );
  OAI22_X1 U2007 ( .A1(n9281), .A2(n9692), .B1(n8847), .B2(n9697), .ZN(n3674)
         );
  OAI22_X1 U2008 ( .A1(n9278), .A2(n9692), .B1(n8848), .B2(n9697), .ZN(n3658)
         );
  OAI22_X1 U2009 ( .A1(n9275), .A2(n9692), .B1(n8849), .B2(n9697), .ZN(n3642)
         );
  OAI22_X1 U2010 ( .A1(n9272), .A2(n9691), .B1(n8850), .B2(n9698), .ZN(n3626)
         );
  OAI22_X1 U2011 ( .A1(n9269), .A2(n9691), .B1(n8851), .B2(n9698), .ZN(n3610)
         );
  OAI22_X1 U2012 ( .A1(n9266), .A2(n9691), .B1(n8852), .B2(n9698), .ZN(n3594)
         );
  OAI22_X1 U2013 ( .A1(n9263), .A2(n9691), .B1(n8853), .B2(n9698), .ZN(n3578)
         );
  OAI22_X1 U2014 ( .A1(n9260), .A2(n9691), .B1(n8854), .B2(n9699), .ZN(n3562)
         );
  OAI22_X1 U2015 ( .A1(n9257), .A2(n9691), .B1(n8855), .B2(n9699), .ZN(n3546)
         );
  OAI22_X1 U2016 ( .A1(n9254), .A2(n9691), .B1(n8856), .B2(n9699), .ZN(n3530)
         );
  OAI22_X1 U2017 ( .A1(n9251), .A2(n9691), .B1(n8857), .B2(n9699), .ZN(n3514)
         );
  OAI22_X1 U2018 ( .A1(n9248), .A2(n9691), .B1(n8858), .B2(n9700), .ZN(n3498)
         );
  OAI22_X1 U2019 ( .A1(n9245), .A2(n9691), .B1(n8859), .B2(n9700), .ZN(n3482)
         );
  OAI22_X1 U2020 ( .A1(n9242), .A2(n9691), .B1(n8860), .B2(n9700), .ZN(n3466)
         );
  OAI22_X1 U2021 ( .A1(n9239), .A2(n9691), .B1(n8861), .B2(n9700), .ZN(n3450)
         );
  OAI22_X1 U2022 ( .A1(n9332), .A2(n9681), .B1(n8918), .B2(n9682), .ZN(n3944)
         );
  OAI22_X1 U2023 ( .A1(n9329), .A2(n9680), .B1(n8919), .B2(n9682), .ZN(n3928)
         );
  OAI22_X1 U2024 ( .A1(n9326), .A2(n9681), .B1(n8920), .B2(n9682), .ZN(n3912)
         );
  OAI22_X1 U2025 ( .A1(n9323), .A2(n9680), .B1(n8921), .B2(n9682), .ZN(n3896)
         );
  OAI22_X1 U2026 ( .A1(n9320), .A2(n9681), .B1(n8922), .B2(n9683), .ZN(n3880)
         );
  OAI22_X1 U2027 ( .A1(n9317), .A2(n9680), .B1(n8923), .B2(n9683), .ZN(n3864)
         );
  OAI22_X1 U2028 ( .A1(n9314), .A2(n9681), .B1(n8924), .B2(n9683), .ZN(n3848)
         );
  OAI22_X1 U2029 ( .A1(n9311), .A2(n9680), .B1(n8925), .B2(n9683), .ZN(n3832)
         );
  OAI22_X1 U2030 ( .A1(n9308), .A2(n9681), .B1(n8926), .B2(n9684), .ZN(n3816)
         );
  OAI22_X1 U2031 ( .A1(n9305), .A2(n9681), .B1(n8927), .B2(n9684), .ZN(n3800)
         );
  OAI22_X1 U2032 ( .A1(n9302), .A2(n9681), .B1(n8928), .B2(n9684), .ZN(n3784)
         );
  OAI22_X1 U2033 ( .A1(n9299), .A2(n9681), .B1(n8929), .B2(n9684), .ZN(n3768)
         );
  OAI22_X1 U2034 ( .A1(n9296), .A2(n9681), .B1(n8930), .B2(n9685), .ZN(n3752)
         );
  OAI22_X1 U2035 ( .A1(n9293), .A2(n9681), .B1(n8931), .B2(n9685), .ZN(n3736)
         );
  OAI22_X1 U2036 ( .A1(n9290), .A2(n9681), .B1(n8932), .B2(n9685), .ZN(n3720)
         );
  OAI22_X1 U2037 ( .A1(n9287), .A2(n9681), .B1(n8933), .B2(n9685), .ZN(n3704)
         );
  OAI22_X1 U2038 ( .A1(n9284), .A2(n9681), .B1(n8934), .B2(n9686), .ZN(n3688)
         );
  OAI22_X1 U2039 ( .A1(n9281), .A2(n9681), .B1(n8935), .B2(n9686), .ZN(n3672)
         );
  OAI22_X1 U2040 ( .A1(n9278), .A2(n9681), .B1(n8936), .B2(n9686), .ZN(n3656)
         );
  OAI22_X1 U2041 ( .A1(n9275), .A2(n9681), .B1(n8937), .B2(n9686), .ZN(n3640)
         );
  OAI22_X1 U2042 ( .A1(n9272), .A2(n9680), .B1(n8938), .B2(n9687), .ZN(n3624)
         );
  OAI22_X1 U2043 ( .A1(n9269), .A2(n9680), .B1(n8939), .B2(n9687), .ZN(n3608)
         );
  OAI22_X1 U2044 ( .A1(n9266), .A2(n9680), .B1(n8940), .B2(n9687), .ZN(n3592)
         );
  OAI22_X1 U2045 ( .A1(n9263), .A2(n9680), .B1(n8941), .B2(n9687), .ZN(n3576)
         );
  OAI22_X1 U2046 ( .A1(n9260), .A2(n9680), .B1(n8942), .B2(n9688), .ZN(n3560)
         );
  OAI22_X1 U2047 ( .A1(n9257), .A2(n9680), .B1(n8943), .B2(n9688), .ZN(n3544)
         );
  OAI22_X1 U2048 ( .A1(n9254), .A2(n9680), .B1(n8944), .B2(n9688), .ZN(n3528)
         );
  OAI22_X1 U2049 ( .A1(n9251), .A2(n9680), .B1(n8945), .B2(n9688), .ZN(n3512)
         );
  OAI22_X1 U2050 ( .A1(n9248), .A2(n9680), .B1(n8946), .B2(n9689), .ZN(n3496)
         );
  OAI22_X1 U2051 ( .A1(n9245), .A2(n9680), .B1(n8947), .B2(n9689), .ZN(n3480)
         );
  OAI22_X1 U2052 ( .A1(n9242), .A2(n9680), .B1(n8948), .B2(n9689), .ZN(n3464)
         );
  OAI22_X1 U2053 ( .A1(n9239), .A2(n9680), .B1(n8949), .B2(n9689), .ZN(n3448)
         );
  OAI22_X1 U2054 ( .A1(n9875), .A2(n9331), .B1(n2349), .B2(n9867), .ZN(n9174)
         );
  OAI22_X1 U2055 ( .A1(n9875), .A2(n9328), .B1(n2341), .B2(n9867), .ZN(n9175)
         );
  OAI22_X1 U2056 ( .A1(n9874), .A2(n9325), .B1(n2333), .B2(n9867), .ZN(n9176)
         );
  OAI22_X1 U2057 ( .A1(n9874), .A2(n9322), .B1(n2325), .B2(n9867), .ZN(n9177)
         );
  OAI22_X1 U2058 ( .A1(n9874), .A2(n9319), .B1(n2317), .B2(n9867), .ZN(n9178)
         );
  OAI22_X1 U2059 ( .A1(n9874), .A2(n9316), .B1(n2309), .B2(n9867), .ZN(n9179)
         );
  OAI22_X1 U2060 ( .A1(n9874), .A2(n9313), .B1(n2301), .B2(n9867), .ZN(n9180)
         );
  OAI22_X1 U2061 ( .A1(n9873), .A2(n9310), .B1(n2293), .B2(n9867), .ZN(n9181)
         );
  OAI22_X1 U2062 ( .A1(n9873), .A2(n9307), .B1(n2285), .B2(n9867), .ZN(n9182)
         );
  OAI22_X1 U2063 ( .A1(n9873), .A2(n9304), .B1(n2277), .B2(n9867), .ZN(n9183)
         );
  OAI22_X1 U2064 ( .A1(n9873), .A2(n9301), .B1(n2269), .B2(n9867), .ZN(n9184)
         );
  OAI22_X1 U2065 ( .A1(n9873), .A2(n9298), .B1(n2261), .B2(n9867), .ZN(n9185)
         );
  OAI22_X1 U2066 ( .A1(n9872), .A2(n9295), .B1(n2253), .B2(n9868), .ZN(n9186)
         );
  OAI22_X1 U2067 ( .A1(n9872), .A2(n9292), .B1(n2245), .B2(n9868), .ZN(n9187)
         );
  OAI22_X1 U2068 ( .A1(n9872), .A2(n9289), .B1(n2237), .B2(n9868), .ZN(n9188)
         );
  OAI22_X1 U2069 ( .A1(n9872), .A2(n9286), .B1(n2229), .B2(n9868), .ZN(n9189)
         );
  OAI22_X1 U2070 ( .A1(n9872), .A2(n9283), .B1(n2221), .B2(n9868), .ZN(n9190)
         );
  OAI22_X1 U2071 ( .A1(n9871), .A2(n9280), .B1(n2213), .B2(n9868), .ZN(n9191)
         );
  OAI22_X1 U2072 ( .A1(n9871), .A2(n9277), .B1(n2205), .B2(n9868), .ZN(n9192)
         );
  OAI22_X1 U2073 ( .A1(n9871), .A2(n9274), .B1(n2197), .B2(n9868), .ZN(n9193)
         );
  OAI22_X1 U2074 ( .A1(n9871), .A2(n9271), .B1(n2189), .B2(n9868), .ZN(n9194)
         );
  OAI22_X1 U2075 ( .A1(n9871), .A2(n9268), .B1(n2181), .B2(n9868), .ZN(n9195)
         );
  OAI22_X1 U2076 ( .A1(n9870), .A2(n9265), .B1(n2173), .B2(n9868), .ZN(n9196)
         );
  OAI22_X1 U2077 ( .A1(n9870), .A2(n9262), .B1(n2165), .B2(n9868), .ZN(n9197)
         );
  OAI22_X1 U2078 ( .A1(n9312), .A2(n9548), .B1(n8246), .B2(n9556), .ZN(n3045)
         );
  OAI22_X1 U2079 ( .A1(n9309), .A2(n9548), .B1(n8247), .B2(n9555), .ZN(n3046)
         );
  OAI22_X1 U2080 ( .A1(n9306), .A2(n9548), .B1(n8248), .B2(n9555), .ZN(n3047)
         );
  OAI22_X1 U2081 ( .A1(n9303), .A2(n9548), .B1(n8249), .B2(n9555), .ZN(n3048)
         );
  OAI22_X1 U2082 ( .A1(n9300), .A2(n9548), .B1(n8250), .B2(n9555), .ZN(n3049)
         );
  OAI22_X1 U2083 ( .A1(n9297), .A2(n9549), .B1(n8251), .B2(n9554), .ZN(n3050)
         );
  OAI22_X1 U2084 ( .A1(n9294), .A2(n9549), .B1(n8252), .B2(n9554), .ZN(n3051)
         );
  OAI22_X1 U2085 ( .A1(n9291), .A2(n9549), .B1(n8253), .B2(n9554), .ZN(n3052)
         );
  OAI22_X1 U2086 ( .A1(n9288), .A2(n9549), .B1(n8254), .B2(n9554), .ZN(n3053)
         );
  OAI22_X1 U2087 ( .A1(n9285), .A2(n9549), .B1(n8255), .B2(n9553), .ZN(n3054)
         );
  OAI22_X1 U2088 ( .A1(n9282), .A2(n9549), .B1(n8256), .B2(n9553), .ZN(n3055)
         );
  OAI22_X1 U2089 ( .A1(n9279), .A2(n9549), .B1(n8257), .B2(n9553), .ZN(n3056)
         );
  OAI22_X1 U2090 ( .A1(n9276), .A2(n9549), .B1(n8258), .B2(n9553), .ZN(n3057)
         );
  OAI22_X1 U2091 ( .A1(n9273), .A2(n9549), .B1(n8259), .B2(n9552), .ZN(n3058)
         );
  OAI22_X1 U2092 ( .A1(n9270), .A2(n9549), .B1(n8260), .B2(n9552), .ZN(n3059)
         );
  OAI22_X1 U2093 ( .A1(n9267), .A2(n9549), .B1(n8261), .B2(n9552), .ZN(n3060)
         );
  OAI22_X1 U2094 ( .A1(n9264), .A2(n9549), .B1(n8262), .B2(n9552), .ZN(n3061)
         );
  OAI22_X1 U2095 ( .A1(n9260), .A2(n9636), .B1(n8311), .B2(n9639), .ZN(n3318)
         );
  OAI22_X1 U2096 ( .A1(n9257), .A2(n9637), .B1(n8312), .B2(n9639), .ZN(n3319)
         );
  OAI22_X1 U2097 ( .A1(n9254), .A2(n9636), .B1(n8313), .B2(n9639), .ZN(n3320)
         );
  OAI22_X1 U2098 ( .A1(n9251), .A2(n9637), .B1(n8314), .B2(n9639), .ZN(n3321)
         );
  OAI22_X1 U2099 ( .A1(n9248), .A2(n9636), .B1(n8315), .B2(n9638), .ZN(n3322)
         );
  OAI22_X1 U2100 ( .A1(n9245), .A2(n9637), .B1(n8316), .B2(n9638), .ZN(n3323)
         );
  OAI22_X1 U2101 ( .A1(n9242), .A2(n9636), .B1(n8317), .B2(n9638), .ZN(n3324)
         );
  OAI22_X1 U2102 ( .A1(n9239), .A2(n9637), .B1(n8318), .B2(n9638), .ZN(n3325)
         );
  OAI22_X1 U2103 ( .A1(n9261), .A2(n9549), .B1(n8327), .B2(n9551), .ZN(n3062)
         );
  OAI22_X1 U2104 ( .A1(n9258), .A2(n9548), .B1(n8328), .B2(n9551), .ZN(n3063)
         );
  OAI22_X1 U2105 ( .A1(n9255), .A2(n9549), .B1(n8329), .B2(n9551), .ZN(n3064)
         );
  OAI22_X1 U2106 ( .A1(n9252), .A2(n9548), .B1(n8330), .B2(n9551), .ZN(n3065)
         );
  OAI22_X1 U2107 ( .A1(n9249), .A2(n9549), .B1(n8331), .B2(n9550), .ZN(n3066)
         );
  OAI22_X1 U2108 ( .A1(n9246), .A2(n9548), .B1(n8332), .B2(n9550), .ZN(n3067)
         );
  OAI22_X1 U2109 ( .A1(n9243), .A2(n9549), .B1(n8333), .B2(n9550), .ZN(n3068)
         );
  OAI22_X1 U2110 ( .A1(n9240), .A2(n9548), .B1(n8334), .B2(n9550), .ZN(n3069)
         );
  OAI22_X1 U2111 ( .A1(n9331), .A2(n9769), .B1(n8375), .B2(n9770), .ZN(n3957)
         );
  OAI22_X1 U2112 ( .A1(n9328), .A2(n9768), .B1(n8376), .B2(n9770), .ZN(n3941)
         );
  OAI22_X1 U2113 ( .A1(n9325), .A2(n9769), .B1(n8377), .B2(n9770), .ZN(n3925)
         );
  OAI22_X1 U2114 ( .A1(n9322), .A2(n9768), .B1(n8378), .B2(n9770), .ZN(n3909)
         );
  OAI22_X1 U2115 ( .A1(n9319), .A2(n9769), .B1(n8379), .B2(n9771), .ZN(n3893)
         );
  OAI22_X1 U2116 ( .A1(n9316), .A2(n9768), .B1(n8380), .B2(n9771), .ZN(n3877)
         );
  OAI22_X1 U2117 ( .A1(n9313), .A2(n9769), .B1(n8381), .B2(n9771), .ZN(n3861)
         );
  OAI22_X1 U2118 ( .A1(n9310), .A2(n9768), .B1(n8382), .B2(n9771), .ZN(n3845)
         );
  OAI22_X1 U2119 ( .A1(n9307), .A2(n9769), .B1(n8383), .B2(n9772), .ZN(n3829)
         );
  OAI22_X1 U2120 ( .A1(n9304), .A2(n9769), .B1(n8384), .B2(n9772), .ZN(n3813)
         );
  OAI22_X1 U2121 ( .A1(n9301), .A2(n9769), .B1(n8385), .B2(n9772), .ZN(n3797)
         );
  OAI22_X1 U2122 ( .A1(n9298), .A2(n9769), .B1(n8386), .B2(n9772), .ZN(n3781)
         );
  OAI22_X1 U2123 ( .A1(n9295), .A2(n9769), .B1(n8387), .B2(n9773), .ZN(n3765)
         );
  OAI22_X1 U2124 ( .A1(n9292), .A2(n9769), .B1(n8388), .B2(n9773), .ZN(n3749)
         );
  OAI22_X1 U2125 ( .A1(n9289), .A2(n9769), .B1(n8389), .B2(n9773), .ZN(n3733)
         );
  OAI22_X1 U2126 ( .A1(n9286), .A2(n9769), .B1(n8390), .B2(n9773), .ZN(n3717)
         );
  OAI22_X1 U2127 ( .A1(n9283), .A2(n9769), .B1(n8391), .B2(n9774), .ZN(n3701)
         );
  OAI22_X1 U2128 ( .A1(n9280), .A2(n9769), .B1(n8392), .B2(n9774), .ZN(n3685)
         );
  OAI22_X1 U2129 ( .A1(n9277), .A2(n9769), .B1(n8393), .B2(n9774), .ZN(n3669)
         );
  OAI22_X1 U2130 ( .A1(n9274), .A2(n9769), .B1(n8394), .B2(n9774), .ZN(n3653)
         );
  OAI22_X1 U2131 ( .A1(n9271), .A2(n9768), .B1(n8395), .B2(n9775), .ZN(n3637)
         );
  OAI22_X1 U2132 ( .A1(n9268), .A2(n9768), .B1(n8396), .B2(n9775), .ZN(n3621)
         );
  OAI22_X1 U2133 ( .A1(n9265), .A2(n9768), .B1(n8397), .B2(n9775), .ZN(n3605)
         );
  OAI22_X1 U2134 ( .A1(n9262), .A2(n9768), .B1(n8398), .B2(n9775), .ZN(n3589)
         );
  OAI22_X1 U2135 ( .A1(n9259), .A2(n9768), .B1(n8399), .B2(n9776), .ZN(n3573)
         );
  OAI22_X1 U2136 ( .A1(n9256), .A2(n9768), .B1(n8400), .B2(n9776), .ZN(n3557)
         );
  OAI22_X1 U2137 ( .A1(n9253), .A2(n9768), .B1(n8401), .B2(n9776), .ZN(n3541)
         );
  OAI22_X1 U2138 ( .A1(n9250), .A2(n9768), .B1(n8402), .B2(n9776), .ZN(n3525)
         );
  OAI22_X1 U2139 ( .A1(n9247), .A2(n9768), .B1(n8403), .B2(n9777), .ZN(n3509)
         );
  OAI22_X1 U2140 ( .A1(n9244), .A2(n9768), .B1(n8404), .B2(n9777), .ZN(n3493)
         );
  OAI22_X1 U2141 ( .A1(n9241), .A2(n9768), .B1(n8405), .B2(n9777), .ZN(n3477)
         );
  OAI22_X1 U2142 ( .A1(n9238), .A2(n9768), .B1(n8406), .B2(n9777), .ZN(n3461)
         );
  OAI22_X1 U2143 ( .A1(n9333), .A2(n9548), .B1(n8471), .B2(n9557), .ZN(n3038)
         );
  OAI22_X1 U2144 ( .A1(n9330), .A2(n9548), .B1(n8472), .B2(n9557), .ZN(n3039)
         );
  OAI22_X1 U2145 ( .A1(n9327), .A2(n9548), .B1(n8473), .B2(n9557), .ZN(n3040)
         );
  OAI22_X1 U2146 ( .A1(n9324), .A2(n9548), .B1(n8474), .B2(n9557), .ZN(n3041)
         );
  OAI22_X1 U2147 ( .A1(n9321), .A2(n9548), .B1(n8475), .B2(n9556), .ZN(n3042)
         );
  OAI22_X1 U2148 ( .A1(n9318), .A2(n9548), .B1(n8476), .B2(n9556), .ZN(n3043)
         );
  OAI22_X1 U2149 ( .A1(n9315), .A2(n9548), .B1(n8477), .B2(n9556), .ZN(n3044)
         );
  OAI22_X1 U2150 ( .A1(n9333), .A2(n9559), .B1(n8478), .B2(n9568), .ZN(n3070)
         );
  OAI22_X1 U2151 ( .A1(n9330), .A2(n9559), .B1(n8479), .B2(n9568), .ZN(n3071)
         );
  OAI22_X1 U2152 ( .A1(n9327), .A2(n9559), .B1(n8480), .B2(n9568), .ZN(n3072)
         );
  OAI22_X1 U2153 ( .A1(n9324), .A2(n9559), .B1(n8481), .B2(n9568), .ZN(n3073)
         );
  OAI22_X1 U2154 ( .A1(n9321), .A2(n9559), .B1(n8482), .B2(n9567), .ZN(n3074)
         );
  OAI22_X1 U2155 ( .A1(n9318), .A2(n9559), .B1(n8483), .B2(n9567), .ZN(n3075)
         );
  OAI22_X1 U2156 ( .A1(n9315), .A2(n9559), .B1(n8484), .B2(n9567), .ZN(n3076)
         );
  OAI22_X1 U2157 ( .A1(n9312), .A2(n9559), .B1(n8485), .B2(n9567), .ZN(n3077)
         );
  OAI22_X1 U2158 ( .A1(n9309), .A2(n9559), .B1(n8486), .B2(n9566), .ZN(n3078)
         );
  OAI22_X1 U2159 ( .A1(n9306), .A2(n9559), .B1(n8487), .B2(n9566), .ZN(n3079)
         );
  OAI22_X1 U2160 ( .A1(n9303), .A2(n9559), .B1(n8488), .B2(n9566), .ZN(n3080)
         );
  OAI22_X1 U2161 ( .A1(n9300), .A2(n9559), .B1(n8489), .B2(n9566), .ZN(n3081)
         );
  OAI22_X1 U2162 ( .A1(n9297), .A2(n9560), .B1(n8490), .B2(n9565), .ZN(n3082)
         );
  OAI22_X1 U2163 ( .A1(n9294), .A2(n9560), .B1(n8491), .B2(n9565), .ZN(n3083)
         );
  OAI22_X1 U2164 ( .A1(n9291), .A2(n9560), .B1(n8492), .B2(n9565), .ZN(n3084)
         );
  OAI22_X1 U2165 ( .A1(n9288), .A2(n9560), .B1(n8493), .B2(n9565), .ZN(n3085)
         );
  OAI22_X1 U2166 ( .A1(n9285), .A2(n9560), .B1(n8494), .B2(n9564), .ZN(n3086)
         );
  OAI22_X1 U2167 ( .A1(n9282), .A2(n9560), .B1(n8495), .B2(n9564), .ZN(n3087)
         );
  OAI22_X1 U2168 ( .A1(n9279), .A2(n9560), .B1(n8496), .B2(n9564), .ZN(n3088)
         );
  OAI22_X1 U2169 ( .A1(n9276), .A2(n9560), .B1(n8497), .B2(n9564), .ZN(n3089)
         );
  OAI22_X1 U2170 ( .A1(n9273), .A2(n9560), .B1(n8498), .B2(n9563), .ZN(n3090)
         );
  OAI22_X1 U2171 ( .A1(n9270), .A2(n9560), .B1(n8499), .B2(n9563), .ZN(n3091)
         );
  OAI22_X1 U2172 ( .A1(n9267), .A2(n9560), .B1(n8500), .B2(n9563), .ZN(n3092)
         );
  OAI22_X1 U2173 ( .A1(n9264), .A2(n9560), .B1(n8501), .B2(n9563), .ZN(n3093)
         );
  OAI22_X1 U2174 ( .A1(n9261), .A2(n9559), .B1(n8502), .B2(n9562), .ZN(n3094)
         );
  OAI22_X1 U2175 ( .A1(n9258), .A2(n9560), .B1(n8503), .B2(n9562), .ZN(n3095)
         );
  OAI22_X1 U2176 ( .A1(n9255), .A2(n9559), .B1(n8504), .B2(n9562), .ZN(n3096)
         );
  OAI22_X1 U2177 ( .A1(n9252), .A2(n9560), .B1(n8505), .B2(n9562), .ZN(n3097)
         );
  OAI22_X1 U2178 ( .A1(n9249), .A2(n9559), .B1(n8506), .B2(n9561), .ZN(n3098)
         );
  OAI22_X1 U2179 ( .A1(n9246), .A2(n9560), .B1(n8507), .B2(n9561), .ZN(n3099)
         );
  OAI22_X1 U2180 ( .A1(n9243), .A2(n9559), .B1(n8508), .B2(n9561), .ZN(n3100)
         );
  OAI22_X1 U2181 ( .A1(n9240), .A2(n9560), .B1(n8509), .B2(n9561), .ZN(n3101)
         );
  OAI22_X1 U2182 ( .A1(n9330), .A2(n9581), .B1(n8567), .B2(n9590), .ZN(n3135)
         );
  OAI22_X1 U2183 ( .A1(n9327), .A2(n9581), .B1(n8568), .B2(n9590), .ZN(n3136)
         );
  OAI22_X1 U2184 ( .A1(n9324), .A2(n9581), .B1(n8569), .B2(n9590), .ZN(n3137)
         );
  OAI22_X1 U2185 ( .A1(n9321), .A2(n9581), .B1(n8570), .B2(n9589), .ZN(n3138)
         );
  OAI22_X1 U2186 ( .A1(n9318), .A2(n9581), .B1(n8571), .B2(n9589), .ZN(n3139)
         );
  OAI22_X1 U2187 ( .A1(n9315), .A2(n9581), .B1(n8572), .B2(n9589), .ZN(n3140)
         );
  OAI22_X1 U2188 ( .A1(n9312), .A2(n9581), .B1(n8573), .B2(n9589), .ZN(n3141)
         );
  OAI22_X1 U2189 ( .A1(n9309), .A2(n9581), .B1(n8574), .B2(n9588), .ZN(n3142)
         );
  OAI22_X1 U2190 ( .A1(n9306), .A2(n9581), .B1(n8575), .B2(n9588), .ZN(n3143)
         );
  OAI22_X1 U2191 ( .A1(n9303), .A2(n9581), .B1(n8576), .B2(n9588), .ZN(n3144)
         );
  OAI22_X1 U2192 ( .A1(n9300), .A2(n9581), .B1(n8577), .B2(n9588), .ZN(n3145)
         );
  OAI22_X1 U2193 ( .A1(n9297), .A2(n9582), .B1(n8578), .B2(n9587), .ZN(n3146)
         );
  OAI22_X1 U2194 ( .A1(n9294), .A2(n9582), .B1(n8579), .B2(n9587), .ZN(n3147)
         );
  OAI22_X1 U2195 ( .A1(n9291), .A2(n9582), .B1(n8580), .B2(n9587), .ZN(n3148)
         );
  OAI22_X1 U2196 ( .A1(n9288), .A2(n9582), .B1(n8581), .B2(n9587), .ZN(n3149)
         );
  OAI22_X1 U2197 ( .A1(n9285), .A2(n9582), .B1(n8582), .B2(n9586), .ZN(n3150)
         );
  OAI22_X1 U2198 ( .A1(n9282), .A2(n9582), .B1(n8583), .B2(n9586), .ZN(n3151)
         );
  OAI22_X1 U2199 ( .A1(n9279), .A2(n9582), .B1(n8584), .B2(n9586), .ZN(n3152)
         );
  OAI22_X1 U2200 ( .A1(n9276), .A2(n9582), .B1(n8585), .B2(n9586), .ZN(n3153)
         );
  OAI22_X1 U2201 ( .A1(n9273), .A2(n9582), .B1(n8586), .B2(n9585), .ZN(n3154)
         );
  OAI22_X1 U2202 ( .A1(n9270), .A2(n9582), .B1(n8587), .B2(n9585), .ZN(n3155)
         );
  OAI22_X1 U2203 ( .A1(n9267), .A2(n9582), .B1(n8588), .B2(n9585), .ZN(n3156)
         );
  OAI22_X1 U2204 ( .A1(n9264), .A2(n9582), .B1(n8589), .B2(n9585), .ZN(n3157)
         );
  OAI22_X1 U2205 ( .A1(n9261), .A2(n9581), .B1(n8590), .B2(n9584), .ZN(n3158)
         );
  OAI22_X1 U2206 ( .A1(n9258), .A2(n9582), .B1(n8591), .B2(n9584), .ZN(n3159)
         );
  OAI22_X1 U2207 ( .A1(n9255), .A2(n9581), .B1(n8592), .B2(n9584), .ZN(n3160)
         );
  OAI22_X1 U2208 ( .A1(n9252), .A2(n9582), .B1(n8593), .B2(n9584), .ZN(n3161)
         );
  OAI22_X1 U2209 ( .A1(n9249), .A2(n9581), .B1(n8594), .B2(n9583), .ZN(n3162)
         );
  OAI22_X1 U2210 ( .A1(n9246), .A2(n9582), .B1(n8595), .B2(n9583), .ZN(n3163)
         );
  OAI22_X1 U2211 ( .A1(n9243), .A2(n9581), .B1(n8596), .B2(n9583), .ZN(n3164)
         );
  OAI22_X1 U2212 ( .A1(n9240), .A2(n9582), .B1(n8597), .B2(n9583), .ZN(n3165)
         );
  OAI22_X1 U2213 ( .A1(n9329), .A2(n9636), .B1(n8775), .B2(n9645), .ZN(n3295)
         );
  OAI22_X1 U2214 ( .A1(n9326), .A2(n9636), .B1(n8776), .B2(n9645), .ZN(n3296)
         );
  OAI22_X1 U2215 ( .A1(n9323), .A2(n9636), .B1(n8777), .B2(n9645), .ZN(n3297)
         );
  OAI22_X1 U2216 ( .A1(n9320), .A2(n9636), .B1(n8778), .B2(n9644), .ZN(n3298)
         );
  OAI22_X1 U2217 ( .A1(n9317), .A2(n9636), .B1(n8779), .B2(n9644), .ZN(n3299)
         );
  OAI22_X1 U2218 ( .A1(n9311), .A2(n9636), .B1(n8781), .B2(n9644), .ZN(n3301)
         );
  OAI22_X1 U2219 ( .A1(n9308), .A2(n9636), .B1(n8782), .B2(n9643), .ZN(n3302)
         );
  OAI22_X1 U2220 ( .A1(n9305), .A2(n9636), .B1(n8783), .B2(n9643), .ZN(n3303)
         );
  OAI22_X1 U2221 ( .A1(n9302), .A2(n9636), .B1(n8784), .B2(n9643), .ZN(n3304)
         );
  OAI22_X1 U2222 ( .A1(n9299), .A2(n9636), .B1(n8785), .B2(n9643), .ZN(n3305)
         );
  OAI22_X1 U2223 ( .A1(n9296), .A2(n9637), .B1(n8786), .B2(n9642), .ZN(n3306)
         );
  OAI22_X1 U2224 ( .A1(n9290), .A2(n9637), .B1(n8788), .B2(n9642), .ZN(n3308)
         );
  OAI22_X1 U2225 ( .A1(n9287), .A2(n9637), .B1(n8789), .B2(n9642), .ZN(n3309)
         );
  OAI22_X1 U2226 ( .A1(n9284), .A2(n9637), .B1(n8790), .B2(n9641), .ZN(n3310)
         );
  OAI22_X1 U2227 ( .A1(n9278), .A2(n9637), .B1(n8792), .B2(n9641), .ZN(n3312)
         );
  OAI22_X1 U2228 ( .A1(n9275), .A2(n9637), .B1(n8793), .B2(n9641), .ZN(n3313)
         );
  OAI22_X1 U2229 ( .A1(n9272), .A2(n9637), .B1(n8794), .B2(n9640), .ZN(n3314)
         );
  OAI22_X1 U2230 ( .A1(n9269), .A2(n9637), .B1(n8795), .B2(n9640), .ZN(n3315)
         );
  OAI22_X1 U2231 ( .A1(n9266), .A2(n9637), .B1(n8796), .B2(n9640), .ZN(n3316)
         );
  OAI22_X1 U2232 ( .A1(n9263), .A2(n9637), .B1(n8797), .B2(n9640), .ZN(n3317)
         );
  OAI22_X1 U2233 ( .A1(n9332), .A2(n9647), .B1(n8798), .B2(n9656), .ZN(n3326)
         );
  OAI22_X1 U2234 ( .A1(n9329), .A2(n9647), .B1(n8799), .B2(n9656), .ZN(n3327)
         );
  OAI22_X1 U2235 ( .A1(n9326), .A2(n9647), .B1(n8800), .B2(n9656), .ZN(n3328)
         );
  OAI22_X1 U2236 ( .A1(n9323), .A2(n9647), .B1(n8801), .B2(n9656), .ZN(n3329)
         );
  OAI22_X1 U2237 ( .A1(n9320), .A2(n9647), .B1(n8802), .B2(n9655), .ZN(n3330)
         );
  OAI22_X1 U2238 ( .A1(n9317), .A2(n9647), .B1(n8803), .B2(n9655), .ZN(n3331)
         );
  OAI22_X1 U2239 ( .A1(n9314), .A2(n9647), .B1(n8804), .B2(n9655), .ZN(n3332)
         );
  OAI22_X1 U2240 ( .A1(n9311), .A2(n9647), .B1(n8805), .B2(n9655), .ZN(n3333)
         );
  OAI22_X1 U2241 ( .A1(n9308), .A2(n9647), .B1(n8806), .B2(n9654), .ZN(n3334)
         );
  OAI22_X1 U2242 ( .A1(n9305), .A2(n9647), .B1(n8807), .B2(n9654), .ZN(n3335)
         );
  OAI22_X1 U2243 ( .A1(n9302), .A2(n9647), .B1(n8808), .B2(n9654), .ZN(n3336)
         );
  OAI22_X1 U2244 ( .A1(n9299), .A2(n9647), .B1(n8809), .B2(n9654), .ZN(n3337)
         );
  OAI22_X1 U2245 ( .A1(n9296), .A2(n9648), .B1(n8810), .B2(n9653), .ZN(n3338)
         );
  OAI22_X1 U2246 ( .A1(n9293), .A2(n9648), .B1(n8811), .B2(n9653), .ZN(n3339)
         );
  OAI22_X1 U2247 ( .A1(n9290), .A2(n9648), .B1(n8812), .B2(n9653), .ZN(n3340)
         );
  OAI22_X1 U2248 ( .A1(n9287), .A2(n9648), .B1(n8813), .B2(n9653), .ZN(n3341)
         );
  OAI22_X1 U2249 ( .A1(n9284), .A2(n9648), .B1(n8814), .B2(n9652), .ZN(n3342)
         );
  OAI22_X1 U2250 ( .A1(n9281), .A2(n9648), .B1(n8815), .B2(n9652), .ZN(n3343)
         );
  OAI22_X1 U2251 ( .A1(n9278), .A2(n9648), .B1(n8816), .B2(n9652), .ZN(n3344)
         );
  OAI22_X1 U2252 ( .A1(n9275), .A2(n9648), .B1(n8817), .B2(n9652), .ZN(n3345)
         );
  OAI22_X1 U2253 ( .A1(n9272), .A2(n9648), .B1(n8818), .B2(n9651), .ZN(n3346)
         );
  OAI22_X1 U2254 ( .A1(n9269), .A2(n9648), .B1(n8819), .B2(n9651), .ZN(n3347)
         );
  OAI22_X1 U2255 ( .A1(n9266), .A2(n9648), .B1(n8820), .B2(n9651), .ZN(n3348)
         );
  OAI22_X1 U2256 ( .A1(n9263), .A2(n9648), .B1(n8821), .B2(n9651), .ZN(n3349)
         );
  OAI22_X1 U2257 ( .A1(n9260), .A2(n9647), .B1(n8822), .B2(n9650), .ZN(n3350)
         );
  OAI22_X1 U2258 ( .A1(n9257), .A2(n9648), .B1(n8823), .B2(n9650), .ZN(n3351)
         );
  OAI22_X1 U2259 ( .A1(n9254), .A2(n9647), .B1(n8824), .B2(n9650), .ZN(n3352)
         );
  OAI22_X1 U2260 ( .A1(n9251), .A2(n9648), .B1(n8825), .B2(n9650), .ZN(n3353)
         );
  OAI22_X1 U2261 ( .A1(n9248), .A2(n9647), .B1(n8826), .B2(n9649), .ZN(n3354)
         );
  OAI22_X1 U2262 ( .A1(n9245), .A2(n9648), .B1(n8827), .B2(n9649), .ZN(n3355)
         );
  OAI22_X1 U2263 ( .A1(n9242), .A2(n9647), .B1(n8828), .B2(n9649), .ZN(n3356)
         );
  OAI22_X1 U2264 ( .A1(n9239), .A2(n9648), .B1(n8829), .B2(n9649), .ZN(n3357)
         );
  OAI22_X1 U2265 ( .A1(n9332), .A2(n9669), .B1(n8886), .B2(n9678), .ZN(n3390)
         );
  OAI22_X1 U2266 ( .A1(n9329), .A2(n9669), .B1(n8887), .B2(n9678), .ZN(n3391)
         );
  OAI22_X1 U2267 ( .A1(n9326), .A2(n9669), .B1(n8888), .B2(n9678), .ZN(n3392)
         );
  OAI22_X1 U2268 ( .A1(n9323), .A2(n9669), .B1(n8889), .B2(n9678), .ZN(n3393)
         );
  OAI22_X1 U2269 ( .A1(n9320), .A2(n9669), .B1(n8890), .B2(n9677), .ZN(n3394)
         );
  OAI22_X1 U2270 ( .A1(n9317), .A2(n9669), .B1(n8891), .B2(n9677), .ZN(n3395)
         );
  OAI22_X1 U2271 ( .A1(n9314), .A2(n9669), .B1(n8892), .B2(n9677), .ZN(n3396)
         );
  OAI22_X1 U2272 ( .A1(n9311), .A2(n9669), .B1(n8893), .B2(n9677), .ZN(n3397)
         );
  OAI22_X1 U2273 ( .A1(n9308), .A2(n9669), .B1(n8894), .B2(n9676), .ZN(n3398)
         );
  OAI22_X1 U2274 ( .A1(n9305), .A2(n9669), .B1(n8895), .B2(n9676), .ZN(n3399)
         );
  OAI22_X1 U2275 ( .A1(n9302), .A2(n9669), .B1(n8896), .B2(n9676), .ZN(n3400)
         );
  OAI22_X1 U2276 ( .A1(n9299), .A2(n9669), .B1(n8897), .B2(n9676), .ZN(n3401)
         );
  OAI22_X1 U2277 ( .A1(n9296), .A2(n9670), .B1(n8898), .B2(n9675), .ZN(n3402)
         );
  OAI22_X1 U2278 ( .A1(n9293), .A2(n9670), .B1(n8899), .B2(n9675), .ZN(n3403)
         );
  OAI22_X1 U2279 ( .A1(n9290), .A2(n9670), .B1(n8900), .B2(n9675), .ZN(n3404)
         );
  OAI22_X1 U2280 ( .A1(n9287), .A2(n9670), .B1(n8901), .B2(n9675), .ZN(n3405)
         );
  OAI22_X1 U2281 ( .A1(n9284), .A2(n9670), .B1(n8902), .B2(n9674), .ZN(n3406)
         );
  OAI22_X1 U2282 ( .A1(n9281), .A2(n9670), .B1(n8903), .B2(n9674), .ZN(n3407)
         );
  OAI22_X1 U2283 ( .A1(n9278), .A2(n9670), .B1(n8904), .B2(n9674), .ZN(n3408)
         );
  OAI22_X1 U2284 ( .A1(n9275), .A2(n9670), .B1(n8905), .B2(n9674), .ZN(n3409)
         );
  OAI22_X1 U2285 ( .A1(n9272), .A2(n9670), .B1(n8906), .B2(n9673), .ZN(n3410)
         );
  OAI22_X1 U2286 ( .A1(n9269), .A2(n9670), .B1(n8907), .B2(n9673), .ZN(n3411)
         );
  OAI22_X1 U2287 ( .A1(n9266), .A2(n9670), .B1(n8908), .B2(n9673), .ZN(n3412)
         );
  OAI22_X1 U2288 ( .A1(n9263), .A2(n9670), .B1(n8909), .B2(n9673), .ZN(n3413)
         );
  OAI22_X1 U2289 ( .A1(n9260), .A2(n9669), .B1(n8910), .B2(n9672), .ZN(n3414)
         );
  OAI22_X1 U2290 ( .A1(n9257), .A2(n9670), .B1(n8911), .B2(n9672), .ZN(n3415)
         );
  OAI22_X1 U2291 ( .A1(n9254), .A2(n9669), .B1(n8912), .B2(n9672), .ZN(n3416)
         );
  OAI22_X1 U2292 ( .A1(n9251), .A2(n9670), .B1(n8913), .B2(n9672), .ZN(n3417)
         );
  OAI22_X1 U2293 ( .A1(n9248), .A2(n9669), .B1(n8914), .B2(n9671), .ZN(n3418)
         );
  OAI22_X1 U2294 ( .A1(n9245), .A2(n9670), .B1(n8915), .B2(n9671), .ZN(n3419)
         );
  OAI22_X1 U2295 ( .A1(n9242), .A2(n9669), .B1(n8916), .B2(n9671), .ZN(n3420)
         );
  OAI22_X1 U2296 ( .A1(n9239), .A2(n9670), .B1(n8917), .B2(n9671), .ZN(n3421)
         );
  OAI22_X1 U2297 ( .A1(n9331), .A2(n9846), .B1(n8244), .B2(n9847), .ZN(n9141)
         );
  OAI22_X1 U2298 ( .A1(n9328), .A2(n9845), .B1(n8242), .B2(n9847), .ZN(n9140)
         );
  OAI22_X1 U2299 ( .A1(n9325), .A2(n9846), .B1(n8240), .B2(n9847), .ZN(n9139)
         );
  OAI22_X1 U2300 ( .A1(n9322), .A2(n9845), .B1(n8238), .B2(n9847), .ZN(n9138)
         );
  OAI22_X1 U2301 ( .A1(n9319), .A2(n9846), .B1(n8236), .B2(n9848), .ZN(n9137)
         );
  OAI22_X1 U2302 ( .A1(n9316), .A2(n9845), .B1(n8234), .B2(n9848), .ZN(n9136)
         );
  OAI22_X1 U2303 ( .A1(n9313), .A2(n9846), .B1(n8232), .B2(n9848), .ZN(n9135)
         );
  OAI22_X1 U2304 ( .A1(n9310), .A2(n9845), .B1(n8230), .B2(n9848), .ZN(n9134)
         );
  OAI22_X1 U2305 ( .A1(n9307), .A2(n9846), .B1(n8228), .B2(n9849), .ZN(n9133)
         );
  OAI22_X1 U2306 ( .A1(n9304), .A2(n9846), .B1(n8226), .B2(n9849), .ZN(n9132)
         );
  OAI22_X1 U2307 ( .A1(n9301), .A2(n9846), .B1(n8224), .B2(n9849), .ZN(n9131)
         );
  OAI22_X1 U2308 ( .A1(n9298), .A2(n9846), .B1(n8222), .B2(n9849), .ZN(n9130)
         );
  OAI22_X1 U2309 ( .A1(n9295), .A2(n9846), .B1(n8220), .B2(n9850), .ZN(n9129)
         );
  OAI22_X1 U2310 ( .A1(n9292), .A2(n9846), .B1(n8218), .B2(n9850), .ZN(n9128)
         );
  OAI22_X1 U2311 ( .A1(n9289), .A2(n9846), .B1(n8216), .B2(n9850), .ZN(n9127)
         );
  OAI22_X1 U2312 ( .A1(n9286), .A2(n9846), .B1(n8214), .B2(n9850), .ZN(n9126)
         );
  OAI22_X1 U2313 ( .A1(n9283), .A2(n9846), .B1(n8212), .B2(n9851), .ZN(n9125)
         );
  OAI22_X1 U2314 ( .A1(n9280), .A2(n9846), .B1(n8210), .B2(n9851), .ZN(n9124)
         );
  OAI22_X1 U2315 ( .A1(n9277), .A2(n9846), .B1(n8208), .B2(n9851), .ZN(n9123)
         );
  OAI22_X1 U2316 ( .A1(n9274), .A2(n9846), .B1(n8206), .B2(n9851), .ZN(n9122)
         );
  OAI22_X1 U2317 ( .A1(n9271), .A2(n9845), .B1(n8204), .B2(n9852), .ZN(n9121)
         );
  OAI22_X1 U2318 ( .A1(n9268), .A2(n9845), .B1(n8202), .B2(n9852), .ZN(n9120)
         );
  OAI22_X1 U2319 ( .A1(n9265), .A2(n9845), .B1(n8200), .B2(n9852), .ZN(n9119)
         );
  OAI22_X1 U2320 ( .A1(n9262), .A2(n9845), .B1(n8198), .B2(n9852), .ZN(n9118)
         );
  OAI22_X1 U2321 ( .A1(n9260), .A2(n9614), .B1(n8287), .B2(n9617), .ZN(n3254)
         );
  OAI22_X1 U2322 ( .A1(n9257), .A2(n9615), .B1(n8288), .B2(n9617), .ZN(n3255)
         );
  OAI22_X1 U2323 ( .A1(n9254), .A2(n9614), .B1(n8289), .B2(n9617), .ZN(n3256)
         );
  OAI22_X1 U2324 ( .A1(n9251), .A2(n9615), .B1(n8290), .B2(n9617), .ZN(n3257)
         );
  OAI22_X1 U2325 ( .A1(n9248), .A2(n9614), .B1(n8291), .B2(n9616), .ZN(n3258)
         );
  OAI22_X1 U2326 ( .A1(n9245), .A2(n9615), .B1(n8292), .B2(n9616), .ZN(n3259)
         );
  OAI22_X1 U2327 ( .A1(n9242), .A2(n9614), .B1(n8293), .B2(n9616), .ZN(n3260)
         );
  OAI22_X1 U2328 ( .A1(n9239), .A2(n9615), .B1(n8294), .B2(n9616), .ZN(n3261)
         );
  OAI22_X1 U2329 ( .A1(n9260), .A2(n9658), .B1(n8303), .B2(n9661), .ZN(n3382)
         );
  OAI22_X1 U2330 ( .A1(n9257), .A2(n9659), .B1(n8304), .B2(n9661), .ZN(n3383)
         );
  OAI22_X1 U2331 ( .A1(n9254), .A2(n9658), .B1(n8305), .B2(n9661), .ZN(n3384)
         );
  OAI22_X1 U2332 ( .A1(n9251), .A2(n9659), .B1(n8306), .B2(n9661), .ZN(n3385)
         );
  OAI22_X1 U2333 ( .A1(n9248), .A2(n9658), .B1(n8307), .B2(n9660), .ZN(n3386)
         );
  OAI22_X1 U2334 ( .A1(n9245), .A2(n9659), .B1(n8308), .B2(n9660), .ZN(n3387)
         );
  OAI22_X1 U2335 ( .A1(n9242), .A2(n9658), .B1(n8309), .B2(n9660), .ZN(n3388)
         );
  OAI22_X1 U2336 ( .A1(n9239), .A2(n9659), .B1(n8310), .B2(n9660), .ZN(n3389)
         );
  OAI22_X1 U2337 ( .A1(n9261), .A2(n9570), .B1(n8319), .B2(n9573), .ZN(n3126)
         );
  OAI22_X1 U2338 ( .A1(n9258), .A2(n9571), .B1(n8320), .B2(n9573), .ZN(n3127)
         );
  OAI22_X1 U2339 ( .A1(n9255), .A2(n9570), .B1(n8321), .B2(n9573), .ZN(n3128)
         );
  OAI22_X1 U2340 ( .A1(n9252), .A2(n9571), .B1(n8322), .B2(n9573), .ZN(n3129)
         );
  OAI22_X1 U2341 ( .A1(n9249), .A2(n9570), .B1(n8323), .B2(n9572), .ZN(n3130)
         );
  OAI22_X1 U2342 ( .A1(n9246), .A2(n9571), .B1(n8324), .B2(n9572), .ZN(n3131)
         );
  OAI22_X1 U2343 ( .A1(n9243), .A2(n9570), .B1(n8325), .B2(n9572), .ZN(n3132)
         );
  OAI22_X1 U2344 ( .A1(n9240), .A2(n9571), .B1(n8326), .B2(n9572), .ZN(n3133)
         );
  OAI22_X1 U2345 ( .A1(n9259), .A2(n9845), .B1(n8196), .B2(n9853), .ZN(n9117)
         );
  OAI22_X1 U2346 ( .A1(n9256), .A2(n9845), .B1(n8194), .B2(n9853), .ZN(n9116)
         );
  OAI22_X1 U2347 ( .A1(n9253), .A2(n9845), .B1(n8192), .B2(n9853), .ZN(n9115)
         );
  OAI22_X1 U2348 ( .A1(n9250), .A2(n9845), .B1(n8190), .B2(n9853), .ZN(n9114)
         );
  OAI22_X1 U2349 ( .A1(n9247), .A2(n9845), .B1(n8188), .B2(n9854), .ZN(n9113)
         );
  OAI22_X1 U2350 ( .A1(n9244), .A2(n9845), .B1(n8186), .B2(n9854), .ZN(n9112)
         );
  OAI22_X1 U2351 ( .A1(n9241), .A2(n9845), .B1(n8184), .B2(n9854), .ZN(n9111)
         );
  OAI22_X1 U2352 ( .A1(n9238), .A2(n9845), .B1(n8182), .B2(n9854), .ZN(n9110)
         );
  OAI22_X1 U2353 ( .A1(n9331), .A2(n9780), .B1(n8343), .B2(n9781), .ZN(n3958)
         );
  OAI22_X1 U2354 ( .A1(n9328), .A2(n9779), .B1(n8344), .B2(n9781), .ZN(n3942)
         );
  OAI22_X1 U2355 ( .A1(n9325), .A2(n9780), .B1(n8345), .B2(n9781), .ZN(n3926)
         );
  OAI22_X1 U2356 ( .A1(n9322), .A2(n9779), .B1(n8346), .B2(n9781), .ZN(n3910)
         );
  OAI22_X1 U2357 ( .A1(n9319), .A2(n9780), .B1(n8347), .B2(n9782), .ZN(n3894)
         );
  OAI22_X1 U2358 ( .A1(n9316), .A2(n9779), .B1(n8348), .B2(n9782), .ZN(n3878)
         );
  OAI22_X1 U2359 ( .A1(n9313), .A2(n9780), .B1(n8349), .B2(n9782), .ZN(n3862)
         );
  OAI22_X1 U2360 ( .A1(n9310), .A2(n9779), .B1(n8350), .B2(n9782), .ZN(n3846)
         );
  OAI22_X1 U2361 ( .A1(n9307), .A2(n9780), .B1(n8351), .B2(n9783), .ZN(n3830)
         );
  OAI22_X1 U2362 ( .A1(n9304), .A2(n9780), .B1(n8352), .B2(n9783), .ZN(n3814)
         );
  OAI22_X1 U2363 ( .A1(n9301), .A2(n9780), .B1(n8353), .B2(n9783), .ZN(n3798)
         );
  OAI22_X1 U2364 ( .A1(n9298), .A2(n9780), .B1(n8354), .B2(n9783), .ZN(n3782)
         );
  OAI22_X1 U2365 ( .A1(n9295), .A2(n9780), .B1(n8355), .B2(n9784), .ZN(n3766)
         );
  OAI22_X1 U2366 ( .A1(n9292), .A2(n9780), .B1(n8356), .B2(n9784), .ZN(n3750)
         );
  OAI22_X1 U2367 ( .A1(n9289), .A2(n9780), .B1(n8357), .B2(n9784), .ZN(n3734)
         );
  OAI22_X1 U2368 ( .A1(n9286), .A2(n9780), .B1(n8358), .B2(n9784), .ZN(n3718)
         );
  OAI22_X1 U2369 ( .A1(n9283), .A2(n9780), .B1(n8359), .B2(n9785), .ZN(n3702)
         );
  OAI22_X1 U2370 ( .A1(n9280), .A2(n9780), .B1(n8360), .B2(n9785), .ZN(n3686)
         );
  OAI22_X1 U2371 ( .A1(n9277), .A2(n9780), .B1(n8361), .B2(n9785), .ZN(n3670)
         );
  OAI22_X1 U2372 ( .A1(n9274), .A2(n9780), .B1(n8362), .B2(n9785), .ZN(n3654)
         );
  OAI22_X1 U2373 ( .A1(n9271), .A2(n9779), .B1(n8363), .B2(n9786), .ZN(n3638)
         );
  OAI22_X1 U2374 ( .A1(n9268), .A2(n9779), .B1(n8364), .B2(n9786), .ZN(n3622)
         );
  OAI22_X1 U2375 ( .A1(n9265), .A2(n9779), .B1(n8365), .B2(n9786), .ZN(n3606)
         );
  OAI22_X1 U2376 ( .A1(n9262), .A2(n9779), .B1(n8366), .B2(n9786), .ZN(n3590)
         );
  OAI22_X1 U2377 ( .A1(n9259), .A2(n9779), .B1(n8367), .B2(n9787), .ZN(n3574)
         );
  OAI22_X1 U2378 ( .A1(n9256), .A2(n9779), .B1(n8368), .B2(n9787), .ZN(n3558)
         );
  OAI22_X1 U2379 ( .A1(n9253), .A2(n9779), .B1(n8369), .B2(n9787), .ZN(n3542)
         );
  OAI22_X1 U2380 ( .A1(n9250), .A2(n9779), .B1(n8370), .B2(n9787), .ZN(n3526)
         );
  OAI22_X1 U2381 ( .A1(n9247), .A2(n9779), .B1(n8371), .B2(n9788), .ZN(n3510)
         );
  OAI22_X1 U2382 ( .A1(n9244), .A2(n9779), .B1(n8372), .B2(n9788), .ZN(n3494)
         );
  OAI22_X1 U2383 ( .A1(n9241), .A2(n9779), .B1(n8373), .B2(n9788), .ZN(n3478)
         );
  OAI22_X1 U2384 ( .A1(n9238), .A2(n9779), .B1(n8374), .B2(n9788), .ZN(n3462)
         );
  OAI22_X1 U2385 ( .A1(n9331), .A2(n9758), .B1(n8407), .B2(n9759), .ZN(n3956)
         );
  OAI22_X1 U2386 ( .A1(n9328), .A2(n9757), .B1(n8408), .B2(n9759), .ZN(n3940)
         );
  OAI22_X1 U2387 ( .A1(n9325), .A2(n9758), .B1(n8409), .B2(n9759), .ZN(n3924)
         );
  OAI22_X1 U2388 ( .A1(n9322), .A2(n9757), .B1(n8410), .B2(n9759), .ZN(n3908)
         );
  OAI22_X1 U2389 ( .A1(n9319), .A2(n9758), .B1(n8411), .B2(n9760), .ZN(n3892)
         );
  OAI22_X1 U2390 ( .A1(n9316), .A2(n9757), .B1(n8412), .B2(n9760), .ZN(n3876)
         );
  OAI22_X1 U2391 ( .A1(n9313), .A2(n9758), .B1(n8413), .B2(n9760), .ZN(n3860)
         );
  OAI22_X1 U2392 ( .A1(n9310), .A2(n9757), .B1(n8414), .B2(n9760), .ZN(n3844)
         );
  OAI22_X1 U2393 ( .A1(n9307), .A2(n9758), .B1(n8415), .B2(n9761), .ZN(n3828)
         );
  OAI22_X1 U2394 ( .A1(n9304), .A2(n9758), .B1(n8416), .B2(n9761), .ZN(n3812)
         );
  OAI22_X1 U2395 ( .A1(n9301), .A2(n9758), .B1(n8417), .B2(n9761), .ZN(n3796)
         );
  OAI22_X1 U2396 ( .A1(n9298), .A2(n9758), .B1(n8418), .B2(n9761), .ZN(n3780)
         );
  OAI22_X1 U2397 ( .A1(n9295), .A2(n9758), .B1(n8419), .B2(n9762), .ZN(n3764)
         );
  OAI22_X1 U2398 ( .A1(n9292), .A2(n9758), .B1(n8420), .B2(n9762), .ZN(n3748)
         );
  OAI22_X1 U2399 ( .A1(n9289), .A2(n9758), .B1(n8421), .B2(n9762), .ZN(n3732)
         );
  OAI22_X1 U2400 ( .A1(n9286), .A2(n9758), .B1(n8422), .B2(n9762), .ZN(n3716)
         );
  OAI22_X1 U2401 ( .A1(n9283), .A2(n9758), .B1(n8423), .B2(n9763), .ZN(n3700)
         );
  OAI22_X1 U2402 ( .A1(n9280), .A2(n9758), .B1(n8424), .B2(n9763), .ZN(n3684)
         );
  OAI22_X1 U2403 ( .A1(n9277), .A2(n9758), .B1(n8425), .B2(n9763), .ZN(n3668)
         );
  OAI22_X1 U2404 ( .A1(n9274), .A2(n9758), .B1(n8426), .B2(n9763), .ZN(n3652)
         );
  OAI22_X1 U2405 ( .A1(n9271), .A2(n9757), .B1(n8427), .B2(n9764), .ZN(n3636)
         );
  OAI22_X1 U2406 ( .A1(n9268), .A2(n9757), .B1(n8428), .B2(n9764), .ZN(n3620)
         );
  OAI22_X1 U2407 ( .A1(n9265), .A2(n9757), .B1(n8429), .B2(n9764), .ZN(n3604)
         );
  OAI22_X1 U2408 ( .A1(n9262), .A2(n9757), .B1(n8430), .B2(n9764), .ZN(n3588)
         );
  OAI22_X1 U2409 ( .A1(n9259), .A2(n9757), .B1(n8431), .B2(n9765), .ZN(n3572)
         );
  OAI22_X1 U2410 ( .A1(n9256), .A2(n9757), .B1(n8432), .B2(n9765), .ZN(n3556)
         );
  OAI22_X1 U2411 ( .A1(n9253), .A2(n9757), .B1(n8433), .B2(n9765), .ZN(n3540)
         );
  OAI22_X1 U2412 ( .A1(n9250), .A2(n9757), .B1(n8434), .B2(n9765), .ZN(n3524)
         );
  OAI22_X1 U2413 ( .A1(n9247), .A2(n9757), .B1(n8435), .B2(n9766), .ZN(n3508)
         );
  OAI22_X1 U2414 ( .A1(n9244), .A2(n9757), .B1(n8436), .B2(n9766), .ZN(n3492)
         );
  OAI22_X1 U2415 ( .A1(n9241), .A2(n9757), .B1(n8437), .B2(n9766), .ZN(n3476)
         );
  OAI22_X1 U2416 ( .A1(n9238), .A2(n9757), .B1(n8438), .B2(n9766), .ZN(n3460)
         );
  OAI22_X1 U2417 ( .A1(n9333), .A2(n9570), .B1(n8542), .B2(n9579), .ZN(n3102)
         );
  OAI22_X1 U2418 ( .A1(n9330), .A2(n9570), .B1(n8543), .B2(n9579), .ZN(n3103)
         );
  OAI22_X1 U2419 ( .A1(n9327), .A2(n9570), .B1(n8544), .B2(n9579), .ZN(n3104)
         );
  OAI22_X1 U2420 ( .A1(n9324), .A2(n9570), .B1(n8545), .B2(n9579), .ZN(n3105)
         );
  OAI22_X1 U2421 ( .A1(n9321), .A2(n9570), .B1(n8546), .B2(n9578), .ZN(n3106)
         );
  OAI22_X1 U2422 ( .A1(n9318), .A2(n9570), .B1(n8547), .B2(n9578), .ZN(n3107)
         );
  OAI22_X1 U2423 ( .A1(n9315), .A2(n9570), .B1(n8548), .B2(n9578), .ZN(n3108)
         );
  OAI22_X1 U2424 ( .A1(n9312), .A2(n9570), .B1(n8549), .B2(n9578), .ZN(n3109)
         );
  OAI22_X1 U2425 ( .A1(n9309), .A2(n9570), .B1(n8550), .B2(n9577), .ZN(n3110)
         );
  OAI22_X1 U2426 ( .A1(n9306), .A2(n9570), .B1(n8551), .B2(n9577), .ZN(n3111)
         );
  OAI22_X1 U2427 ( .A1(n9303), .A2(n9570), .B1(n8552), .B2(n9577), .ZN(n3112)
         );
  OAI22_X1 U2428 ( .A1(n9300), .A2(n9570), .B1(n8553), .B2(n9577), .ZN(n3113)
         );
  OAI22_X1 U2429 ( .A1(n9297), .A2(n9571), .B1(n8554), .B2(n9576), .ZN(n3114)
         );
  OAI22_X1 U2430 ( .A1(n9294), .A2(n9571), .B1(n8555), .B2(n9576), .ZN(n3115)
         );
  OAI22_X1 U2431 ( .A1(n9291), .A2(n9571), .B1(n8556), .B2(n9576), .ZN(n3116)
         );
  OAI22_X1 U2432 ( .A1(n9288), .A2(n9571), .B1(n8557), .B2(n9576), .ZN(n3117)
         );
  OAI22_X1 U2433 ( .A1(n9285), .A2(n9571), .B1(n8558), .B2(n9575), .ZN(n3118)
         );
  OAI22_X1 U2434 ( .A1(n9282), .A2(n9571), .B1(n8559), .B2(n9575), .ZN(n3119)
         );
  OAI22_X1 U2435 ( .A1(n9279), .A2(n9571), .B1(n8560), .B2(n9575), .ZN(n3120)
         );
  OAI22_X1 U2436 ( .A1(n9276), .A2(n9571), .B1(n8561), .B2(n9575), .ZN(n3121)
         );
  OAI22_X1 U2437 ( .A1(n9273), .A2(n9571), .B1(n8562), .B2(n9574), .ZN(n3122)
         );
  OAI22_X1 U2438 ( .A1(n9270), .A2(n9571), .B1(n8563), .B2(n9574), .ZN(n3123)
         );
  OAI22_X1 U2439 ( .A1(n9267), .A2(n9571), .B1(n8564), .B2(n9574), .ZN(n3124)
         );
  OAI22_X1 U2440 ( .A1(n9264), .A2(n9571), .B1(n8565), .B2(n9574), .ZN(n3125)
         );
  OAI22_X1 U2441 ( .A1(n9332), .A2(n9614), .B1(n8718), .B2(n9623), .ZN(n3230)
         );
  OAI22_X1 U2442 ( .A1(n9329), .A2(n9614), .B1(n8719), .B2(n9623), .ZN(n3231)
         );
  OAI22_X1 U2443 ( .A1(n9326), .A2(n9614), .B1(n8720), .B2(n9623), .ZN(n3232)
         );
  OAI22_X1 U2444 ( .A1(n9323), .A2(n9614), .B1(n8721), .B2(n9623), .ZN(n3233)
         );
  OAI22_X1 U2445 ( .A1(n9320), .A2(n9614), .B1(n8722), .B2(n9622), .ZN(n3234)
         );
  OAI22_X1 U2446 ( .A1(n9317), .A2(n9614), .B1(n8723), .B2(n9622), .ZN(n3235)
         );
  OAI22_X1 U2447 ( .A1(n9314), .A2(n9614), .B1(n8724), .B2(n9622), .ZN(n3236)
         );
  OAI22_X1 U2448 ( .A1(n9311), .A2(n9614), .B1(n8725), .B2(n9622), .ZN(n3237)
         );
  OAI22_X1 U2449 ( .A1(n9308), .A2(n9614), .B1(n8726), .B2(n9621), .ZN(n3238)
         );
  OAI22_X1 U2450 ( .A1(n9305), .A2(n9614), .B1(n8727), .B2(n9621), .ZN(n3239)
         );
  OAI22_X1 U2451 ( .A1(n9302), .A2(n9614), .B1(n8728), .B2(n9621), .ZN(n3240)
         );
  OAI22_X1 U2452 ( .A1(n9299), .A2(n9614), .B1(n8729), .B2(n9621), .ZN(n3241)
         );
  OAI22_X1 U2453 ( .A1(n9296), .A2(n9615), .B1(n8730), .B2(n9620), .ZN(n3242)
         );
  OAI22_X1 U2454 ( .A1(n9293), .A2(n9615), .B1(n8731), .B2(n9620), .ZN(n3243)
         );
  OAI22_X1 U2455 ( .A1(n9290), .A2(n9615), .B1(n8732), .B2(n9620), .ZN(n3244)
         );
  OAI22_X1 U2456 ( .A1(n9287), .A2(n9615), .B1(n8733), .B2(n9620), .ZN(n3245)
         );
  OAI22_X1 U2457 ( .A1(n9284), .A2(n9615), .B1(n8734), .B2(n9619), .ZN(n3246)
         );
  OAI22_X1 U2458 ( .A1(n9281), .A2(n9615), .B1(n8735), .B2(n9619), .ZN(n3247)
         );
  OAI22_X1 U2459 ( .A1(n9278), .A2(n9615), .B1(n8736), .B2(n9619), .ZN(n3248)
         );
  OAI22_X1 U2460 ( .A1(n9275), .A2(n9615), .B1(n8737), .B2(n9619), .ZN(n3249)
         );
  OAI22_X1 U2461 ( .A1(n9272), .A2(n9615), .B1(n8738), .B2(n9618), .ZN(n3250)
         );
  OAI22_X1 U2462 ( .A1(n9269), .A2(n9615), .B1(n8739), .B2(n9618), .ZN(n3251)
         );
  OAI22_X1 U2463 ( .A1(n9266), .A2(n9615), .B1(n8740), .B2(n9618), .ZN(n3252)
         );
  OAI22_X1 U2464 ( .A1(n9263), .A2(n9615), .B1(n8741), .B2(n9618), .ZN(n3253)
         );
  OAI22_X1 U2465 ( .A1(n9328), .A2(n9812), .B1(n8243), .B2(n9821), .ZN(n9015)
         );
  OAI22_X1 U2466 ( .A1(n9325), .A2(n9812), .B1(n8241), .B2(n9821), .ZN(n9016)
         );
  OAI22_X1 U2467 ( .A1(n9322), .A2(n9812), .B1(n8239), .B2(n9821), .ZN(n9017)
         );
  OAI22_X1 U2468 ( .A1(n9319), .A2(n9812), .B1(n8237), .B2(n9820), .ZN(n9018)
         );
  OAI22_X1 U2469 ( .A1(n9316), .A2(n9812), .B1(n8235), .B2(n9820), .ZN(n9019)
         );
  OAI22_X1 U2470 ( .A1(n9310), .A2(n9812), .B1(n8231), .B2(n9820), .ZN(n9021)
         );
  OAI22_X1 U2471 ( .A1(n9307), .A2(n9812), .B1(n8229), .B2(n9819), .ZN(n9022)
         );
  OAI22_X1 U2472 ( .A1(n9304), .A2(n9812), .B1(n8227), .B2(n9819), .ZN(n9023)
         );
  OAI22_X1 U2473 ( .A1(n9301), .A2(n9812), .B1(n8225), .B2(n9819), .ZN(n9024)
         );
  OAI22_X1 U2474 ( .A1(n9298), .A2(n9812), .B1(n8223), .B2(n9819), .ZN(n9025)
         );
  OAI22_X1 U2475 ( .A1(n9295), .A2(n9813), .B1(n8221), .B2(n9818), .ZN(n9026)
         );
  OAI22_X1 U2476 ( .A1(n9289), .A2(n9813), .B1(n8217), .B2(n9818), .ZN(n9028)
         );
  OAI22_X1 U2477 ( .A1(n9286), .A2(n9813), .B1(n8215), .B2(n9818), .ZN(n9029)
         );
  OAI22_X1 U2478 ( .A1(n9283), .A2(n9813), .B1(n8213), .B2(n9817), .ZN(n9030)
         );
  OAI22_X1 U2479 ( .A1(n9277), .A2(n9813), .B1(n8209), .B2(n9817), .ZN(n9032)
         );
  OAI22_X1 U2480 ( .A1(n9274), .A2(n9813), .B1(n8207), .B2(n9817), .ZN(n9033)
         );
  OAI22_X1 U2481 ( .A1(n9271), .A2(n9813), .B1(n8205), .B2(n9816), .ZN(n9034)
         );
  OAI22_X1 U2482 ( .A1(n9268), .A2(n9813), .B1(n8203), .B2(n9816), .ZN(n9035)
         );
  OAI22_X1 U2483 ( .A1(n9265), .A2(n9813), .B1(n8201), .B2(n9816), .ZN(n9036)
         );
  OAI22_X1 U2484 ( .A1(n9262), .A2(n9813), .B1(n8199), .B2(n9816), .ZN(n9037)
         );
  OAI22_X1 U2485 ( .A1(n9259), .A2(n9812), .B1(n8197), .B2(n9815), .ZN(n9038)
         );
  OAI22_X1 U2486 ( .A1(n9256), .A2(n9813), .B1(n8195), .B2(n9815), .ZN(n9039)
         );
  OAI22_X1 U2487 ( .A1(n9253), .A2(n9812), .B1(n8193), .B2(n9815), .ZN(n9040)
         );
  OAI22_X1 U2488 ( .A1(n9250), .A2(n9813), .B1(n8191), .B2(n9815), .ZN(n9041)
         );
  OAI22_X1 U2489 ( .A1(n9247), .A2(n9812), .B1(n8189), .B2(n9814), .ZN(n9042)
         );
  OAI22_X1 U2490 ( .A1(n9244), .A2(n9813), .B1(n8187), .B2(n9814), .ZN(n9043)
         );
  OAI22_X1 U2491 ( .A1(n9241), .A2(n9812), .B1(n8185), .B2(n9814), .ZN(n9044)
         );
  OAI22_X1 U2492 ( .A1(n9238), .A2(n9813), .B1(n8183), .B2(n9814), .ZN(n9045)
         );
  OAI22_X1 U2493 ( .A1(n9332), .A2(n9658), .B1(n8862), .B2(n9667), .ZN(n3358)
         );
  OAI22_X1 U2494 ( .A1(n9329), .A2(n9658), .B1(n8863), .B2(n9667), .ZN(n3359)
         );
  OAI22_X1 U2495 ( .A1(n9326), .A2(n9658), .B1(n8864), .B2(n9667), .ZN(n3360)
         );
  OAI22_X1 U2496 ( .A1(n9323), .A2(n9658), .B1(n8865), .B2(n9667), .ZN(n3361)
         );
  OAI22_X1 U2497 ( .A1(n9320), .A2(n9658), .B1(n8866), .B2(n9666), .ZN(n3362)
         );
  OAI22_X1 U2498 ( .A1(n9317), .A2(n9658), .B1(n8867), .B2(n9666), .ZN(n3363)
         );
  OAI22_X1 U2499 ( .A1(n9314), .A2(n9658), .B1(n8868), .B2(n9666), .ZN(n3364)
         );
  OAI22_X1 U2500 ( .A1(n9311), .A2(n9658), .B1(n8869), .B2(n9666), .ZN(n3365)
         );
  OAI22_X1 U2501 ( .A1(n9308), .A2(n9658), .B1(n8870), .B2(n9665), .ZN(n3366)
         );
  OAI22_X1 U2502 ( .A1(n9305), .A2(n9658), .B1(n8871), .B2(n9665), .ZN(n3367)
         );
  OAI22_X1 U2503 ( .A1(n9302), .A2(n9658), .B1(n8872), .B2(n9665), .ZN(n3368)
         );
  OAI22_X1 U2504 ( .A1(n9299), .A2(n9658), .B1(n8873), .B2(n9665), .ZN(n3369)
         );
  OAI22_X1 U2505 ( .A1(n9296), .A2(n9659), .B1(n8874), .B2(n9664), .ZN(n3370)
         );
  OAI22_X1 U2506 ( .A1(n9293), .A2(n9659), .B1(n8875), .B2(n9664), .ZN(n3371)
         );
  OAI22_X1 U2507 ( .A1(n9290), .A2(n9659), .B1(n8876), .B2(n9664), .ZN(n3372)
         );
  OAI22_X1 U2508 ( .A1(n9287), .A2(n9659), .B1(n8877), .B2(n9664), .ZN(n3373)
         );
  OAI22_X1 U2509 ( .A1(n9284), .A2(n9659), .B1(n8878), .B2(n9663), .ZN(n3374)
         );
  OAI22_X1 U2510 ( .A1(n9281), .A2(n9659), .B1(n8879), .B2(n9663), .ZN(n3375)
         );
  OAI22_X1 U2511 ( .A1(n9278), .A2(n9659), .B1(n8880), .B2(n9663), .ZN(n3376)
         );
  OAI22_X1 U2512 ( .A1(n9275), .A2(n9659), .B1(n8881), .B2(n9663), .ZN(n3377)
         );
  OAI22_X1 U2513 ( .A1(n9272), .A2(n9659), .B1(n8882), .B2(n9662), .ZN(n3378)
         );
  OAI22_X1 U2514 ( .A1(n9269), .A2(n9659), .B1(n8883), .B2(n9662), .ZN(n3379)
         );
  OAI22_X1 U2515 ( .A1(n9266), .A2(n9659), .B1(n8884), .B2(n9662), .ZN(n3380)
         );
  OAI22_X1 U2516 ( .A1(n9263), .A2(n9659), .B1(n8885), .B2(n9662), .ZN(n3381)
         );
  OAI22_X1 U2517 ( .A1(n9260), .A2(n9592), .B1(n8295), .B2(n9595), .ZN(n3190)
         );
  OAI22_X1 U2518 ( .A1(n9257), .A2(n9593), .B1(n8296), .B2(n9595), .ZN(n3191)
         );
  OAI22_X1 U2519 ( .A1(n9254), .A2(n9592), .B1(n8297), .B2(n9595), .ZN(n3192)
         );
  OAI22_X1 U2520 ( .A1(n9251), .A2(n9593), .B1(n8298), .B2(n9595), .ZN(n3193)
         );
  OAI22_X1 U2521 ( .A1(n9248), .A2(n9592), .B1(n8299), .B2(n9594), .ZN(n3194)
         );
  OAI22_X1 U2522 ( .A1(n9245), .A2(n9593), .B1(n8300), .B2(n9594), .ZN(n3195)
         );
  OAI22_X1 U2523 ( .A1(n9242), .A2(n9592), .B1(n8301), .B2(n9594), .ZN(n3196)
         );
  OAI22_X1 U2524 ( .A1(n9239), .A2(n9593), .B1(n8302), .B2(n9594), .ZN(n3197)
         );
  OAI22_X1 U2525 ( .A1(n9329), .A2(n9592), .B1(n8631), .B2(n9601), .ZN(n3167)
         );
  OAI22_X1 U2526 ( .A1(n9326), .A2(n9592), .B1(n8632), .B2(n9601), .ZN(n3168)
         );
  OAI22_X1 U2527 ( .A1(n9323), .A2(n9592), .B1(n8633), .B2(n9601), .ZN(n3169)
         );
  OAI22_X1 U2528 ( .A1(n9320), .A2(n9592), .B1(n8634), .B2(n9600), .ZN(n3170)
         );
  OAI22_X1 U2529 ( .A1(n9317), .A2(n9592), .B1(n8635), .B2(n9600), .ZN(n3171)
         );
  OAI22_X1 U2530 ( .A1(n9311), .A2(n9592), .B1(n8637), .B2(n9600), .ZN(n3173)
         );
  OAI22_X1 U2531 ( .A1(n9308), .A2(n9592), .B1(n8638), .B2(n9599), .ZN(n3174)
         );
  OAI22_X1 U2532 ( .A1(n9305), .A2(n9592), .B1(n8639), .B2(n9599), .ZN(n3175)
         );
  OAI22_X1 U2533 ( .A1(n9302), .A2(n9592), .B1(n8640), .B2(n9599), .ZN(n3176)
         );
  OAI22_X1 U2534 ( .A1(n9299), .A2(n9592), .B1(n8641), .B2(n9599), .ZN(n3177)
         );
  OAI22_X1 U2535 ( .A1(n9296), .A2(n9593), .B1(n8642), .B2(n9598), .ZN(n3178)
         );
  OAI22_X1 U2536 ( .A1(n9290), .A2(n9593), .B1(n8644), .B2(n9598), .ZN(n3180)
         );
  OAI22_X1 U2537 ( .A1(n9287), .A2(n9593), .B1(n8645), .B2(n9598), .ZN(n3181)
         );
  OAI22_X1 U2538 ( .A1(n9284), .A2(n9593), .B1(n8646), .B2(n9597), .ZN(n3182)
         );
  OAI22_X1 U2539 ( .A1(n9278), .A2(n9593), .B1(n8648), .B2(n9597), .ZN(n3184)
         );
  OAI22_X1 U2540 ( .A1(n9275), .A2(n9593), .B1(n8649), .B2(n9597), .ZN(n3185)
         );
  OAI22_X1 U2541 ( .A1(n9272), .A2(n9593), .B1(n8650), .B2(n9596), .ZN(n3186)
         );
  OAI22_X1 U2542 ( .A1(n9269), .A2(n9593), .B1(n8651), .B2(n9596), .ZN(n3187)
         );
  OAI22_X1 U2543 ( .A1(n9266), .A2(n9593), .B1(n8652), .B2(n9596), .ZN(n3188)
         );
  OAI22_X1 U2544 ( .A1(n9263), .A2(n9593), .B1(n8653), .B2(n9596), .ZN(n3189)
         );
  OAI22_X1 U2545 ( .A1(n9332), .A2(n9603), .B1(n8654), .B2(n9612), .ZN(n3198)
         );
  OAI22_X1 U2546 ( .A1(n9314), .A2(n9603), .B1(n8660), .B2(n9611), .ZN(n3204)
         );
  OAI22_X1 U2547 ( .A1(n9293), .A2(n9604), .B1(n8667), .B2(n9609), .ZN(n3211)
         );
  OAI22_X1 U2548 ( .A1(n9281), .A2(n9604), .B1(n8671), .B2(n9608), .ZN(n3215)
         );
  OAI22_X1 U2549 ( .A1(n9333), .A2(n9581), .B1(n8566), .B2(n9590), .ZN(n3134)
         );
  OAI22_X1 U2550 ( .A1(n9332), .A2(n9724), .B1(n8598), .B2(n9726), .ZN(n3952)
         );
  OAI22_X1 U2551 ( .A1(n9331), .A2(n9812), .B1(n8245), .B2(n9821), .ZN(n9014)
         );
  OAI22_X1 U2552 ( .A1(n9313), .A2(n9812), .B1(n8233), .B2(n9820), .ZN(n9020)
         );
  OAI22_X1 U2553 ( .A1(n9292), .A2(n9813), .B1(n8219), .B2(n9818), .ZN(n9027)
         );
  OAI22_X1 U2554 ( .A1(n9280), .A2(n9813), .B1(n8211), .B2(n9817), .ZN(n9031)
         );
  OAI22_X1 U2555 ( .A1(n9332), .A2(n9636), .B1(n8774), .B2(n9645), .ZN(n3294)
         );
  OAI22_X1 U2556 ( .A1(n9314), .A2(n9636), .B1(n8780), .B2(n9644), .ZN(n3300)
         );
  OAI22_X1 U2557 ( .A1(n9293), .A2(n9637), .B1(n8787), .B2(n9642), .ZN(n3307)
         );
  OAI22_X1 U2558 ( .A1(n9281), .A2(n9637), .B1(n8791), .B2(n9641), .ZN(n3311)
         );
  OAI22_X1 U2559 ( .A1(n9332), .A2(n9592), .B1(n8630), .B2(n9601), .ZN(n3166)
         );
  OAI22_X1 U2560 ( .A1(n9314), .A2(n9592), .B1(n8636), .B2(n9600), .ZN(n3172)
         );
  OAI22_X1 U2561 ( .A1(n9293), .A2(n9593), .B1(n8643), .B2(n9598), .ZN(n3179)
         );
  OAI22_X1 U2562 ( .A1(n9281), .A2(n9593), .B1(n8647), .B2(n9597), .ZN(n3183)
         );
  OAI22_X1 U2563 ( .A1(n9333), .A2(n9526), .B1(n8263), .B2(n9535), .ZN(n2942)
         );
  OAI22_X1 U2564 ( .A1(n9330), .A2(n9526), .B1(n8264), .B2(n9535), .ZN(n2943)
         );
  OAI22_X1 U2565 ( .A1(n9327), .A2(n9526), .B1(n8265), .B2(n9535), .ZN(n2944)
         );
  OAI22_X1 U2566 ( .A1(n9324), .A2(n9526), .B1(n8266), .B2(n9535), .ZN(n2945)
         );
  OAI22_X1 U2567 ( .A1(n9321), .A2(n9526), .B1(n8267), .B2(n9534), .ZN(n2946)
         );
  OAI22_X1 U2568 ( .A1(n9318), .A2(n9526), .B1(n8268), .B2(n9534), .ZN(n2947)
         );
  OAI22_X1 U2569 ( .A1(n9315), .A2(n9526), .B1(n8269), .B2(n9534), .ZN(n2948)
         );
  OAI22_X1 U2570 ( .A1(n9312), .A2(n9526), .B1(n8270), .B2(n9534), .ZN(n2949)
         );
  OAI22_X1 U2571 ( .A1(n9309), .A2(n9526), .B1(n8271), .B2(n9533), .ZN(n2950)
         );
  OAI22_X1 U2572 ( .A1(n9306), .A2(n9526), .B1(n8272), .B2(n9533), .ZN(n2951)
         );
  OAI22_X1 U2573 ( .A1(n9303), .A2(n9526), .B1(n8273), .B2(n9533), .ZN(n2952)
         );
  OAI22_X1 U2574 ( .A1(n9300), .A2(n9526), .B1(n8274), .B2(n9533), .ZN(n2953)
         );
  OAI22_X1 U2575 ( .A1(n9297), .A2(n9527), .B1(n8275), .B2(n9532), .ZN(n2954)
         );
  OAI22_X1 U2576 ( .A1(n9294), .A2(n9527), .B1(n8276), .B2(n9532), .ZN(n2955)
         );
  OAI22_X1 U2577 ( .A1(n9291), .A2(n9527), .B1(n8277), .B2(n9532), .ZN(n2956)
         );
  OAI22_X1 U2578 ( .A1(n9288), .A2(n9527), .B1(n8278), .B2(n9532), .ZN(n2957)
         );
  OAI22_X1 U2579 ( .A1(n9285), .A2(n9527), .B1(n8279), .B2(n9531), .ZN(n2958)
         );
  OAI22_X1 U2580 ( .A1(n9282), .A2(n9527), .B1(n8280), .B2(n9531), .ZN(n2959)
         );
  OAI22_X1 U2581 ( .A1(n9279), .A2(n9527), .B1(n8281), .B2(n9531), .ZN(n2960)
         );
  OAI22_X1 U2582 ( .A1(n9276), .A2(n9527), .B1(n8282), .B2(n9531), .ZN(n2961)
         );
  OAI22_X1 U2583 ( .A1(n9273), .A2(n9527), .B1(n8283), .B2(n9530), .ZN(n2962)
         );
  OAI22_X1 U2584 ( .A1(n9270), .A2(n9527), .B1(n8284), .B2(n9530), .ZN(n2963)
         );
  OAI22_X1 U2585 ( .A1(n9267), .A2(n9527), .B1(n8285), .B2(n9530), .ZN(n2964)
         );
  OAI22_X1 U2586 ( .A1(n9264), .A2(n9527), .B1(n8286), .B2(n9530), .ZN(n2965)
         );
  OAI22_X1 U2587 ( .A1(n9333), .A2(n9537), .B1(n2350), .B2(n9546), .ZN(n2974)
         );
  OAI22_X1 U2588 ( .A1(n9330), .A2(n9537), .B1(n2342), .B2(n9546), .ZN(n2975)
         );
  OAI22_X1 U2589 ( .A1(n9327), .A2(n9537), .B1(n2334), .B2(n9546), .ZN(n2976)
         );
  OAI22_X1 U2590 ( .A1(n9324), .A2(n9537), .B1(n2326), .B2(n9546), .ZN(n2977)
         );
  OAI22_X1 U2591 ( .A1(n9321), .A2(n9537), .B1(n2318), .B2(n9545), .ZN(n2978)
         );
  OAI22_X1 U2592 ( .A1(n9318), .A2(n9537), .B1(n2310), .B2(n9545), .ZN(n2979)
         );
  OAI22_X1 U2593 ( .A1(n9315), .A2(n9537), .B1(n2302), .B2(n9545), .ZN(n2980)
         );
  OAI22_X1 U2594 ( .A1(n9312), .A2(n9537), .B1(n2294), .B2(n9545), .ZN(n2981)
         );
  OAI22_X1 U2595 ( .A1(n9309), .A2(n9537), .B1(n2286), .B2(n9544), .ZN(n2982)
         );
  OAI22_X1 U2596 ( .A1(n9306), .A2(n9537), .B1(n2278), .B2(n9544), .ZN(n2983)
         );
  OAI22_X1 U2597 ( .A1(n9303), .A2(n9537), .B1(n2270), .B2(n9544), .ZN(n2984)
         );
  OAI22_X1 U2598 ( .A1(n9300), .A2(n9537), .B1(n2262), .B2(n9544), .ZN(n2985)
         );
  OAI22_X1 U2599 ( .A1(n9297), .A2(n9538), .B1(n2254), .B2(n9543), .ZN(n2986)
         );
  OAI22_X1 U2600 ( .A1(n9294), .A2(n9538), .B1(n2246), .B2(n9543), .ZN(n2987)
         );
  OAI22_X1 U2601 ( .A1(n9291), .A2(n9538), .B1(n2238), .B2(n9543), .ZN(n2988)
         );
  OAI22_X1 U2602 ( .A1(n9288), .A2(n9538), .B1(n2230), .B2(n9543), .ZN(n2989)
         );
  OAI22_X1 U2603 ( .A1(n9285), .A2(n9538), .B1(n2222), .B2(n9542), .ZN(n2990)
         );
  OAI22_X1 U2604 ( .A1(n9282), .A2(n9538), .B1(n2214), .B2(n9542), .ZN(n2991)
         );
  OAI22_X1 U2605 ( .A1(n9279), .A2(n9538), .B1(n2206), .B2(n9542), .ZN(n2992)
         );
  OAI22_X1 U2606 ( .A1(n9276), .A2(n9538), .B1(n2198), .B2(n9542), .ZN(n2993)
         );
  OAI22_X1 U2607 ( .A1(n9273), .A2(n9538), .B1(n2190), .B2(n9541), .ZN(n2994)
         );
  OAI22_X1 U2608 ( .A1(n9270), .A2(n9538), .B1(n2182), .B2(n9541), .ZN(n2995)
         );
  OAI22_X1 U2609 ( .A1(n9267), .A2(n9538), .B1(n2174), .B2(n9541), .ZN(n2996)
         );
  OAI22_X1 U2610 ( .A1(n9264), .A2(n9538), .B1(n2166), .B2(n9541), .ZN(n2997)
         );
  OAI22_X1 U2611 ( .A1(n9261), .A2(n9526), .B1(n8335), .B2(n9529), .ZN(n2966)
         );
  OAI22_X1 U2612 ( .A1(n9258), .A2(n9527), .B1(n8336), .B2(n9529), .ZN(n2967)
         );
  OAI22_X1 U2613 ( .A1(n9255), .A2(n9526), .B1(n8337), .B2(n9529), .ZN(n2968)
         );
  OAI22_X1 U2614 ( .A1(n9252), .A2(n9527), .B1(n8338), .B2(n9529), .ZN(n2969)
         );
  OAI22_X1 U2615 ( .A1(n9249), .A2(n9526), .B1(n8339), .B2(n9528), .ZN(n2970)
         );
  OAI22_X1 U2616 ( .A1(n9246), .A2(n9527), .B1(n8340), .B2(n9528), .ZN(n2971)
         );
  OAI22_X1 U2617 ( .A1(n9243), .A2(n9526), .B1(n8341), .B2(n9528), .ZN(n2972)
         );
  OAI22_X1 U2618 ( .A1(n9240), .A2(n9527), .B1(n8342), .B2(n9528), .ZN(n2973)
         );
  OAI22_X1 U2619 ( .A1(n9261), .A2(n9537), .B1(n2158), .B2(n9540), .ZN(n2998)
         );
  OAI22_X1 U2620 ( .A1(n9258), .A2(n9538), .B1(n2150), .B2(n9540), .ZN(n2999)
         );
  OAI22_X1 U2621 ( .A1(n9255), .A2(n9537), .B1(n2142), .B2(n9540), .ZN(n3000)
         );
  OAI22_X1 U2622 ( .A1(n9252), .A2(n9538), .B1(n2134), .B2(n9540), .ZN(n3001)
         );
  OAI22_X1 U2623 ( .A1(n9249), .A2(n9537), .B1(n2126), .B2(n9539), .ZN(n3002)
         );
  OAI22_X1 U2624 ( .A1(n9246), .A2(n9538), .B1(n2118), .B2(n9539), .ZN(n3003)
         );
  OAI22_X1 U2625 ( .A1(n9243), .A2(n9537), .B1(n2110), .B2(n9539), .ZN(n3004)
         );
  OAI22_X1 U2626 ( .A1(n9240), .A2(n9538), .B1(n2102), .B2(n9539), .ZN(n3005)
         );
  OAI22_X1 U2627 ( .A1(n9331), .A2(n9856), .B1(n2348), .B2(n9865), .ZN(n9142)
         );
  OAI22_X1 U2628 ( .A1(n9328), .A2(n9856), .B1(n2340), .B2(n9865), .ZN(n9143)
         );
  OAI22_X1 U2629 ( .A1(n9325), .A2(n9856), .B1(n2332), .B2(n9865), .ZN(n9144)
         );
  OAI22_X1 U2630 ( .A1(n9322), .A2(n9856), .B1(n2324), .B2(n9865), .ZN(n9145)
         );
  OAI22_X1 U2631 ( .A1(n9319), .A2(n9856), .B1(n2316), .B2(n9864), .ZN(n9146)
         );
  OAI22_X1 U2632 ( .A1(n9316), .A2(n9856), .B1(n2308), .B2(n9864), .ZN(n9147)
         );
  OAI22_X1 U2633 ( .A1(n9313), .A2(n9856), .B1(n2300), .B2(n9864), .ZN(n9148)
         );
  OAI22_X1 U2634 ( .A1(n9310), .A2(n9856), .B1(n2292), .B2(n9864), .ZN(n9149)
         );
  OAI22_X1 U2635 ( .A1(n9307), .A2(n9856), .B1(n2284), .B2(n9863), .ZN(n9150)
         );
  OAI22_X1 U2636 ( .A1(n9304), .A2(n9856), .B1(n2276), .B2(n9863), .ZN(n9151)
         );
  OAI22_X1 U2637 ( .A1(n9301), .A2(n9856), .B1(n2268), .B2(n9863), .ZN(n9152)
         );
  OAI22_X1 U2638 ( .A1(n9298), .A2(n9856), .B1(n2260), .B2(n9863), .ZN(n9153)
         );
  OAI22_X1 U2639 ( .A1(n9295), .A2(n9857), .B1(n2252), .B2(n9862), .ZN(n9154)
         );
  OAI22_X1 U2640 ( .A1(n9292), .A2(n9857), .B1(n2244), .B2(n9862), .ZN(n9155)
         );
  OAI22_X1 U2641 ( .A1(n9289), .A2(n9857), .B1(n2236), .B2(n9862), .ZN(n9156)
         );
  OAI22_X1 U2642 ( .A1(n9286), .A2(n9857), .B1(n2228), .B2(n9862), .ZN(n9157)
         );
  OAI22_X1 U2643 ( .A1(n9283), .A2(n9857), .B1(n2220), .B2(n9861), .ZN(n9158)
         );
  OAI22_X1 U2644 ( .A1(n9280), .A2(n9857), .B1(n2212), .B2(n9861), .ZN(n9159)
         );
  OAI22_X1 U2645 ( .A1(n9277), .A2(n9857), .B1(n2204), .B2(n9861), .ZN(n9160)
         );
  OAI22_X1 U2646 ( .A1(n9274), .A2(n9857), .B1(n2196), .B2(n9861), .ZN(n9161)
         );
  OAI22_X1 U2647 ( .A1(n9271), .A2(n9857), .B1(n2188), .B2(n9860), .ZN(n9162)
         );
  OAI22_X1 U2648 ( .A1(n9268), .A2(n9857), .B1(n2180), .B2(n9860), .ZN(n9163)
         );
  OAI22_X1 U2649 ( .A1(n9265), .A2(n9857), .B1(n2172), .B2(n9860), .ZN(n9164)
         );
  OAI22_X1 U2650 ( .A1(n9262), .A2(n9857), .B1(n2164), .B2(n9860), .ZN(n9165)
         );
  OAI22_X1 U2651 ( .A1(n9259), .A2(n9856), .B1(n2156), .B2(n9859), .ZN(n9166)
         );
  OAI22_X1 U2652 ( .A1(n9256), .A2(n9857), .B1(n2148), .B2(n9859), .ZN(n9167)
         );
  OAI22_X1 U2653 ( .A1(n9253), .A2(n9856), .B1(n2140), .B2(n9859), .ZN(n9168)
         );
  OAI22_X1 U2654 ( .A1(n9250), .A2(n9857), .B1(n2132), .B2(n9859), .ZN(n9169)
         );
  OAI22_X1 U2655 ( .A1(n9247), .A2(n9856), .B1(n2124), .B2(n9858), .ZN(n9170)
         );
  OAI22_X1 U2656 ( .A1(n9244), .A2(n9857), .B1(n2116), .B2(n9858), .ZN(n9171)
         );
  OAI22_X1 U2657 ( .A1(n9241), .A2(n9856), .B1(n2108), .B2(n9858), .ZN(n9172)
         );
  OAI22_X1 U2658 ( .A1(n9238), .A2(n9857), .B1(n2100), .B2(n9858), .ZN(n9173)
         );
  OAI22_X1 U2659 ( .A1(n9331), .A2(n9823), .B1(n2355), .B2(n9832), .ZN(n9046)
         );
  OAI22_X1 U2660 ( .A1(n9328), .A2(n9823), .B1(n2347), .B2(n9832), .ZN(n9047)
         );
  OAI22_X1 U2661 ( .A1(n9325), .A2(n9823), .B1(n2339), .B2(n9832), .ZN(n9048)
         );
  OAI22_X1 U2662 ( .A1(n9322), .A2(n9823), .B1(n2331), .B2(n9832), .ZN(n9049)
         );
  OAI22_X1 U2663 ( .A1(n9319), .A2(n9823), .B1(n2323), .B2(n9831), .ZN(n9050)
         );
  OAI22_X1 U2664 ( .A1(n9316), .A2(n9823), .B1(n2315), .B2(n9831), .ZN(n9051)
         );
  OAI22_X1 U2665 ( .A1(n9313), .A2(n9823), .B1(n2307), .B2(n9831), .ZN(n9052)
         );
  OAI22_X1 U2666 ( .A1(n9310), .A2(n9823), .B1(n2299), .B2(n9831), .ZN(n9053)
         );
  OAI22_X1 U2667 ( .A1(n9307), .A2(n9823), .B1(n2291), .B2(n9830), .ZN(n9054)
         );
  OAI22_X1 U2668 ( .A1(n9304), .A2(n9823), .B1(n2283), .B2(n9830), .ZN(n9055)
         );
  OAI22_X1 U2669 ( .A1(n9301), .A2(n9823), .B1(n2275), .B2(n9830), .ZN(n9056)
         );
  OAI22_X1 U2670 ( .A1(n9298), .A2(n9823), .B1(n2267), .B2(n9830), .ZN(n9057)
         );
  OAI22_X1 U2671 ( .A1(n9295), .A2(n9824), .B1(n2259), .B2(n9829), .ZN(n9058)
         );
  OAI22_X1 U2672 ( .A1(n9292), .A2(n9824), .B1(n2251), .B2(n9829), .ZN(n9059)
         );
  OAI22_X1 U2673 ( .A1(n9289), .A2(n9824), .B1(n2243), .B2(n9829), .ZN(n9060)
         );
  OAI22_X1 U2674 ( .A1(n9286), .A2(n9824), .B1(n2235), .B2(n9829), .ZN(n9061)
         );
  OAI22_X1 U2675 ( .A1(n9283), .A2(n9824), .B1(n2227), .B2(n9828), .ZN(n9062)
         );
  OAI22_X1 U2676 ( .A1(n9280), .A2(n9824), .B1(n2219), .B2(n9828), .ZN(n9063)
         );
  OAI22_X1 U2677 ( .A1(n9277), .A2(n9824), .B1(n2211), .B2(n9828), .ZN(n9064)
         );
  OAI22_X1 U2678 ( .A1(n9274), .A2(n9824), .B1(n2203), .B2(n9828), .ZN(n9065)
         );
  OAI22_X1 U2679 ( .A1(n9271), .A2(n9824), .B1(n2195), .B2(n9827), .ZN(n9066)
         );
  OAI22_X1 U2680 ( .A1(n9268), .A2(n9824), .B1(n2187), .B2(n9827), .ZN(n9067)
         );
  OAI22_X1 U2681 ( .A1(n9265), .A2(n9824), .B1(n2179), .B2(n9827), .ZN(n9068)
         );
  OAI22_X1 U2682 ( .A1(n9262), .A2(n9824), .B1(n2171), .B2(n9827), .ZN(n9069)
         );
  OAI22_X1 U2683 ( .A1(n9259), .A2(n9823), .B1(n2163), .B2(n9826), .ZN(n9070)
         );
  OAI22_X1 U2684 ( .A1(n9256), .A2(n9824), .B1(n2155), .B2(n9826), .ZN(n9071)
         );
  OAI22_X1 U2685 ( .A1(n9253), .A2(n9823), .B1(n2147), .B2(n9826), .ZN(n9072)
         );
  OAI22_X1 U2686 ( .A1(n9250), .A2(n9824), .B1(n2139), .B2(n9826), .ZN(n9073)
         );
  OAI22_X1 U2687 ( .A1(n9247), .A2(n9823), .B1(n2131), .B2(n9825), .ZN(n9074)
         );
  OAI22_X1 U2688 ( .A1(n9244), .A2(n9824), .B1(n2123), .B2(n9825), .ZN(n9075)
         );
  OAI22_X1 U2689 ( .A1(n9241), .A2(n9823), .B1(n2115), .B2(n9825), .ZN(n9076)
         );
  OAI22_X1 U2690 ( .A1(n9238), .A2(n9824), .B1(n2107), .B2(n9825), .ZN(n9077)
         );
  OAI22_X1 U2691 ( .A1(n9332), .A2(n9714), .B1(n8686), .B2(n9715), .ZN(n3949)
         );
  OAI22_X1 U2692 ( .A1(n9329), .A2(n9713), .B1(n8687), .B2(n9715), .ZN(n3933)
         );
  OAI22_X1 U2693 ( .A1(n9326), .A2(n9714), .B1(n8688), .B2(n9715), .ZN(n3917)
         );
  OAI22_X1 U2694 ( .A1(n9323), .A2(n9713), .B1(n8689), .B2(n9715), .ZN(n3901)
         );
  OAI22_X1 U2695 ( .A1(n9320), .A2(n9714), .B1(n8690), .B2(n9716), .ZN(n3885)
         );
  OAI22_X1 U2696 ( .A1(n9317), .A2(n9713), .B1(n8691), .B2(n9716), .ZN(n3869)
         );
  OAI22_X1 U2697 ( .A1(n9314), .A2(n9714), .B1(n8692), .B2(n9716), .ZN(n3853)
         );
  OAI22_X1 U2698 ( .A1(n9311), .A2(n9713), .B1(n8693), .B2(n9716), .ZN(n3837)
         );
  OAI22_X1 U2699 ( .A1(n9308), .A2(n9714), .B1(n8694), .B2(n9717), .ZN(n3821)
         );
  OAI22_X1 U2700 ( .A1(n9305), .A2(n9714), .B1(n8695), .B2(n9717), .ZN(n3805)
         );
  OAI22_X1 U2701 ( .A1(n9302), .A2(n9714), .B1(n8696), .B2(n9717), .ZN(n3789)
         );
  OAI22_X1 U2702 ( .A1(n9299), .A2(n9714), .B1(n8697), .B2(n9717), .ZN(n3773)
         );
  OAI22_X1 U2703 ( .A1(n9296), .A2(n9714), .B1(n8698), .B2(n9718), .ZN(n3757)
         );
  OAI22_X1 U2704 ( .A1(n9293), .A2(n9714), .B1(n8699), .B2(n9718), .ZN(n3741)
         );
  OAI22_X1 U2705 ( .A1(n9290), .A2(n9714), .B1(n8700), .B2(n9718), .ZN(n3725)
         );
  OAI22_X1 U2706 ( .A1(n9287), .A2(n9714), .B1(n8701), .B2(n9718), .ZN(n3709)
         );
  OAI22_X1 U2707 ( .A1(n9284), .A2(n9714), .B1(n8702), .B2(n9719), .ZN(n3693)
         );
  OAI22_X1 U2708 ( .A1(n9281), .A2(n9714), .B1(n8703), .B2(n9719), .ZN(n3677)
         );
  OAI22_X1 U2709 ( .A1(n9278), .A2(n9714), .B1(n8704), .B2(n9719), .ZN(n3661)
         );
  OAI22_X1 U2710 ( .A1(n9275), .A2(n9714), .B1(n8705), .B2(n9719), .ZN(n3645)
         );
  OAI22_X1 U2711 ( .A1(n9272), .A2(n9713), .B1(n8706), .B2(n9720), .ZN(n3629)
         );
  OAI22_X1 U2712 ( .A1(n9269), .A2(n9713), .B1(n8707), .B2(n9720), .ZN(n3613)
         );
  OAI22_X1 U2713 ( .A1(n9266), .A2(n9713), .B1(n8708), .B2(n9720), .ZN(n3597)
         );
  OAI22_X1 U2714 ( .A1(n9263), .A2(n9713), .B1(n8709), .B2(n9720), .ZN(n3581)
         );
  OAI22_X1 U2715 ( .A1(n9260), .A2(n9713), .B1(n8710), .B2(n9721), .ZN(n3565)
         );
  OAI22_X1 U2716 ( .A1(n9257), .A2(n9713), .B1(n8711), .B2(n9721), .ZN(n3549)
         );
  OAI22_X1 U2717 ( .A1(n9254), .A2(n9713), .B1(n8712), .B2(n9721), .ZN(n3533)
         );
  OAI22_X1 U2718 ( .A1(n9251), .A2(n9713), .B1(n8713), .B2(n9721), .ZN(n3517)
         );
  OAI22_X1 U2719 ( .A1(n9248), .A2(n9713), .B1(n8714), .B2(n9722), .ZN(n3501)
         );
  OAI22_X1 U2720 ( .A1(n9245), .A2(n9713), .B1(n8715), .B2(n9722), .ZN(n3485)
         );
  OAI22_X1 U2721 ( .A1(n9242), .A2(n9713), .B1(n8716), .B2(n9722), .ZN(n3469)
         );
  OAI22_X1 U2722 ( .A1(n9239), .A2(n9713), .B1(n8717), .B2(n9722), .ZN(n3453)
         );
  OAI22_X1 U2723 ( .A1(n9332), .A2(n9703), .B1(n2354), .B2(n9704), .ZN(n3948)
         );
  OAI22_X1 U2724 ( .A1(n9329), .A2(n9702), .B1(n2346), .B2(n9704), .ZN(n3932)
         );
  OAI22_X1 U2725 ( .A1(n9326), .A2(n9703), .B1(n2338), .B2(n9704), .ZN(n3916)
         );
  OAI22_X1 U2726 ( .A1(n9323), .A2(n9702), .B1(n2330), .B2(n9704), .ZN(n3900)
         );
  OAI22_X1 U2727 ( .A1(n9320), .A2(n9703), .B1(n2322), .B2(n9705), .ZN(n3884)
         );
  OAI22_X1 U2728 ( .A1(n9317), .A2(n9702), .B1(n2314), .B2(n9705), .ZN(n3868)
         );
  OAI22_X1 U2729 ( .A1(n9314), .A2(n9703), .B1(n2306), .B2(n9705), .ZN(n3852)
         );
  OAI22_X1 U2730 ( .A1(n9311), .A2(n9702), .B1(n2298), .B2(n9705), .ZN(n3836)
         );
  OAI22_X1 U2731 ( .A1(n9308), .A2(n9703), .B1(n2290), .B2(n9706), .ZN(n3820)
         );
  OAI22_X1 U2732 ( .A1(n9305), .A2(n9703), .B1(n2282), .B2(n9706), .ZN(n3804)
         );
  OAI22_X1 U2733 ( .A1(n9302), .A2(n9703), .B1(n2274), .B2(n9706), .ZN(n3788)
         );
  OAI22_X1 U2734 ( .A1(n9299), .A2(n9703), .B1(n2266), .B2(n9706), .ZN(n3772)
         );
  OAI22_X1 U2735 ( .A1(n9296), .A2(n9703), .B1(n2258), .B2(n9707), .ZN(n3756)
         );
  OAI22_X1 U2736 ( .A1(n9293), .A2(n9703), .B1(n2250), .B2(n9707), .ZN(n3740)
         );
  OAI22_X1 U2737 ( .A1(n9290), .A2(n9703), .B1(n2242), .B2(n9707), .ZN(n3724)
         );
  OAI22_X1 U2738 ( .A1(n9287), .A2(n9703), .B1(n2234), .B2(n9707), .ZN(n3708)
         );
  OAI22_X1 U2739 ( .A1(n9284), .A2(n9703), .B1(n2226), .B2(n9708), .ZN(n3692)
         );
  OAI22_X1 U2740 ( .A1(n9281), .A2(n9703), .B1(n2218), .B2(n9708), .ZN(n3676)
         );
  OAI22_X1 U2741 ( .A1(n9278), .A2(n9703), .B1(n2210), .B2(n9708), .ZN(n3660)
         );
  OAI22_X1 U2742 ( .A1(n9275), .A2(n9703), .B1(n2202), .B2(n9708), .ZN(n3644)
         );
  OAI22_X1 U2743 ( .A1(n9272), .A2(n9702), .B1(n2194), .B2(n9709), .ZN(n3628)
         );
  OAI22_X1 U2744 ( .A1(n9269), .A2(n9702), .B1(n2186), .B2(n9709), .ZN(n3612)
         );
  OAI22_X1 U2745 ( .A1(n9266), .A2(n9702), .B1(n2178), .B2(n9709), .ZN(n3596)
         );
  OAI22_X1 U2746 ( .A1(n9263), .A2(n9702), .B1(n2170), .B2(n9709), .ZN(n3580)
         );
  OAI22_X1 U2747 ( .A1(n9260), .A2(n9702), .B1(n2162), .B2(n9710), .ZN(n3564)
         );
  OAI22_X1 U2748 ( .A1(n9257), .A2(n9702), .B1(n2154), .B2(n9710), .ZN(n3548)
         );
  OAI22_X1 U2749 ( .A1(n9254), .A2(n9702), .B1(n2146), .B2(n9710), .ZN(n3532)
         );
  OAI22_X1 U2750 ( .A1(n9251), .A2(n9702), .B1(n2138), .B2(n9710), .ZN(n3516)
         );
  OAI22_X1 U2751 ( .A1(n9248), .A2(n9702), .B1(n2130), .B2(n9711), .ZN(n3500)
         );
  OAI22_X1 U2752 ( .A1(n9245), .A2(n9702), .B1(n2122), .B2(n9711), .ZN(n3484)
         );
  OAI22_X1 U2753 ( .A1(n9242), .A2(n9702), .B1(n2114), .B2(n9711), .ZN(n3468)
         );
  OAI22_X1 U2754 ( .A1(n9239), .A2(n9702), .B1(n2106), .B2(n9711), .ZN(n3452)
         );
  OAI22_X1 U2755 ( .A1(n9331), .A2(n9801), .B1(n2353), .B2(n9810), .ZN(n8982)
         );
  OAI22_X1 U2756 ( .A1(n9328), .A2(n9801), .B1(n2345), .B2(n9810), .ZN(n8983)
         );
  OAI22_X1 U2757 ( .A1(n9325), .A2(n9801), .B1(n2337), .B2(n9810), .ZN(n8984)
         );
  OAI22_X1 U2758 ( .A1(n9322), .A2(n9801), .B1(n2329), .B2(n9810), .ZN(n8985)
         );
  OAI22_X1 U2759 ( .A1(n9319), .A2(n9801), .B1(n2321), .B2(n9809), .ZN(n8986)
         );
  OAI22_X1 U2760 ( .A1(n9316), .A2(n9801), .B1(n2313), .B2(n9809), .ZN(n8987)
         );
  OAI22_X1 U2761 ( .A1(n9313), .A2(n9801), .B1(n2305), .B2(n9809), .ZN(n8988)
         );
  OAI22_X1 U2762 ( .A1(n9310), .A2(n9801), .B1(n2297), .B2(n9809), .ZN(n8989)
         );
  OAI22_X1 U2763 ( .A1(n9307), .A2(n9801), .B1(n2289), .B2(n9808), .ZN(n8990)
         );
  OAI22_X1 U2764 ( .A1(n9304), .A2(n9801), .B1(n2281), .B2(n9808), .ZN(n8991)
         );
  OAI22_X1 U2765 ( .A1(n9301), .A2(n9801), .B1(n2273), .B2(n9808), .ZN(n8992)
         );
  OAI22_X1 U2766 ( .A1(n9298), .A2(n9801), .B1(n2265), .B2(n9808), .ZN(n8993)
         );
  OAI22_X1 U2767 ( .A1(n9295), .A2(n9802), .B1(n2257), .B2(n9807), .ZN(n8994)
         );
  OAI22_X1 U2768 ( .A1(n9292), .A2(n9802), .B1(n2249), .B2(n9807), .ZN(n8995)
         );
  OAI22_X1 U2769 ( .A1(n9289), .A2(n9802), .B1(n2241), .B2(n9807), .ZN(n8996)
         );
  OAI22_X1 U2770 ( .A1(n9286), .A2(n9802), .B1(n2233), .B2(n9807), .ZN(n8997)
         );
  OAI22_X1 U2771 ( .A1(n9283), .A2(n9802), .B1(n2225), .B2(n9806), .ZN(n8998)
         );
  OAI22_X1 U2772 ( .A1(n9280), .A2(n9802), .B1(n2217), .B2(n9806), .ZN(n8999)
         );
  OAI22_X1 U2773 ( .A1(n9277), .A2(n9802), .B1(n2209), .B2(n9806), .ZN(n9000)
         );
  OAI22_X1 U2774 ( .A1(n9274), .A2(n9802), .B1(n2201), .B2(n9806), .ZN(n9001)
         );
  OAI22_X1 U2775 ( .A1(n9271), .A2(n9802), .B1(n2193), .B2(n9805), .ZN(n9002)
         );
  OAI22_X1 U2776 ( .A1(n9268), .A2(n9802), .B1(n2185), .B2(n9805), .ZN(n9003)
         );
  OAI22_X1 U2777 ( .A1(n9265), .A2(n9802), .B1(n2177), .B2(n9805), .ZN(n9004)
         );
  OAI22_X1 U2778 ( .A1(n9262), .A2(n9802), .B1(n2169), .B2(n9805), .ZN(n9005)
         );
  OAI22_X1 U2779 ( .A1(n9259), .A2(n9801), .B1(n2161), .B2(n9804), .ZN(n9006)
         );
  OAI22_X1 U2780 ( .A1(n9256), .A2(n9802), .B1(n2153), .B2(n9804), .ZN(n9007)
         );
  OAI22_X1 U2781 ( .A1(n9253), .A2(n9801), .B1(n2145), .B2(n9804), .ZN(n9008)
         );
  OAI22_X1 U2782 ( .A1(n9250), .A2(n9802), .B1(n2137), .B2(n9804), .ZN(n9009)
         );
  OAI22_X1 U2783 ( .A1(n9247), .A2(n9801), .B1(n2129), .B2(n9803), .ZN(n9010)
         );
  OAI22_X1 U2784 ( .A1(n9244), .A2(n9802), .B1(n2121), .B2(n9803), .ZN(n9011)
         );
  OAI22_X1 U2785 ( .A1(n9241), .A2(n9801), .B1(n2113), .B2(n9803), .ZN(n9012)
         );
  OAI22_X1 U2786 ( .A1(n9238), .A2(n9802), .B1(n2105), .B2(n9803), .ZN(n9013)
         );
  OAI22_X1 U2787 ( .A1(n9331), .A2(n9790), .B1(n2352), .B2(n9799), .ZN(n8950)
         );
  OAI22_X1 U2788 ( .A1(n9328), .A2(n9790), .B1(n2344), .B2(n9799), .ZN(n8951)
         );
  OAI22_X1 U2789 ( .A1(n9325), .A2(n9790), .B1(n2336), .B2(n9799), .ZN(n8952)
         );
  OAI22_X1 U2790 ( .A1(n9322), .A2(n9790), .B1(n2328), .B2(n9799), .ZN(n8953)
         );
  OAI22_X1 U2791 ( .A1(n9319), .A2(n9790), .B1(n2320), .B2(n9798), .ZN(n8954)
         );
  OAI22_X1 U2792 ( .A1(n9316), .A2(n9790), .B1(n2312), .B2(n9798), .ZN(n8955)
         );
  OAI22_X1 U2793 ( .A1(n9313), .A2(n9790), .B1(n2304), .B2(n9798), .ZN(n8956)
         );
  OAI22_X1 U2794 ( .A1(n9310), .A2(n9790), .B1(n2296), .B2(n9798), .ZN(n8957)
         );
  OAI22_X1 U2795 ( .A1(n9307), .A2(n9790), .B1(n2288), .B2(n9797), .ZN(n8958)
         );
  OAI22_X1 U2796 ( .A1(n9304), .A2(n9790), .B1(n2280), .B2(n9797), .ZN(n8959)
         );
  OAI22_X1 U2797 ( .A1(n9301), .A2(n9790), .B1(n2272), .B2(n9797), .ZN(n8960)
         );
  OAI22_X1 U2798 ( .A1(n9298), .A2(n9790), .B1(n2264), .B2(n9797), .ZN(n8961)
         );
  OAI22_X1 U2799 ( .A1(n9295), .A2(n9791), .B1(n2256), .B2(n9796), .ZN(n8962)
         );
  OAI22_X1 U2800 ( .A1(n9292), .A2(n9791), .B1(n2248), .B2(n9796), .ZN(n8963)
         );
  OAI22_X1 U2801 ( .A1(n9289), .A2(n9791), .B1(n2240), .B2(n9796), .ZN(n8964)
         );
  OAI22_X1 U2802 ( .A1(n9286), .A2(n9791), .B1(n2232), .B2(n9796), .ZN(n8965)
         );
  OAI22_X1 U2803 ( .A1(n9283), .A2(n9791), .B1(n2224), .B2(n9795), .ZN(n8966)
         );
  OAI22_X1 U2804 ( .A1(n9280), .A2(n9791), .B1(n2216), .B2(n9795), .ZN(n8967)
         );
  OAI22_X1 U2805 ( .A1(n9277), .A2(n9791), .B1(n2208), .B2(n9795), .ZN(n8968)
         );
  OAI22_X1 U2806 ( .A1(n9274), .A2(n9791), .B1(n2200), .B2(n9795), .ZN(n8969)
         );
  OAI22_X1 U2807 ( .A1(n9271), .A2(n9791), .B1(n2192), .B2(n9794), .ZN(n8970)
         );
  OAI22_X1 U2808 ( .A1(n9268), .A2(n9791), .B1(n2184), .B2(n9794), .ZN(n8971)
         );
  OAI22_X1 U2809 ( .A1(n9265), .A2(n9791), .B1(n2176), .B2(n9794), .ZN(n8972)
         );
  OAI22_X1 U2810 ( .A1(n9262), .A2(n9791), .B1(n2168), .B2(n9794), .ZN(n8973)
         );
  OAI22_X1 U2811 ( .A1(n9259), .A2(n9790), .B1(n2160), .B2(n9793), .ZN(n8974)
         );
  OAI22_X1 U2812 ( .A1(n9256), .A2(n9791), .B1(n2152), .B2(n9793), .ZN(n8975)
         );
  OAI22_X1 U2813 ( .A1(n9253), .A2(n9790), .B1(n2144), .B2(n9793), .ZN(n8976)
         );
  OAI22_X1 U2814 ( .A1(n9250), .A2(n9791), .B1(n2136), .B2(n9793), .ZN(n8977)
         );
  OAI22_X1 U2815 ( .A1(n9247), .A2(n9790), .B1(n2128), .B2(n9792), .ZN(n8978)
         );
  OAI22_X1 U2816 ( .A1(n9244), .A2(n9791), .B1(n2120), .B2(n9792), .ZN(n8979)
         );
  OAI22_X1 U2817 ( .A1(n9241), .A2(n9790), .B1(n2112), .B2(n9792), .ZN(n8980)
         );
  OAI22_X1 U2818 ( .A1(n9238), .A2(n9791), .B1(n2104), .B2(n9792), .ZN(n8981)
         );
  NAND2_X1 U2819 ( .A1(n1638), .A2(n1639), .ZN(N1044) );
  NOR4_X1 U2820 ( .A1(n1648), .A2(n1649), .A3(n1650), .A4(n1651), .ZN(n1638)
         );
  NAND2_X1 U2821 ( .A1(n1620), .A2(n1621), .ZN(N1045) );
  NOR4_X1 U2822 ( .A1(n1630), .A2(n1631), .A3(n1632), .A4(n1633), .ZN(n1620)
         );
  NAND2_X1 U2823 ( .A1(n1602), .A2(n1603), .ZN(N1046) );
  NOR4_X1 U2824 ( .A1(n1612), .A2(n1613), .A3(n1614), .A4(n1615), .ZN(n1602)
         );
  NAND2_X1 U2825 ( .A1(n1584), .A2(n1585), .ZN(N1047) );
  NOR4_X1 U2826 ( .A1(n1594), .A2(n1595), .A3(n1596), .A4(n1597), .ZN(n1584)
         );
  NAND2_X1 U2827 ( .A1(n1566), .A2(n1567), .ZN(N1048) );
  NOR4_X1 U2828 ( .A1(n1576), .A2(n1577), .A3(n1578), .A4(n1579), .ZN(n1566)
         );
  NAND2_X1 U2829 ( .A1(n1548), .A2(n1549), .ZN(N1049) );
  NOR4_X1 U2830 ( .A1(n1558), .A2(n1559), .A3(n1560), .A4(n1561), .ZN(n1548)
         );
  NAND2_X1 U2831 ( .A1(n1530), .A2(n1531), .ZN(N1050) );
  NOR4_X1 U2832 ( .A1(n1540), .A2(n1541), .A3(n1542), .A4(n1543), .ZN(n1530)
         );
  NAND2_X1 U2833 ( .A1(n1480), .A2(n1481), .ZN(N1051) );
  NOR4_X1 U2834 ( .A1(n1506), .A2(n1507), .A3(n1508), .A4(n1509), .ZN(n1480)
         );
  NOR4_X1 U2835 ( .A1(n862), .A2(n863), .A3(n864), .A4(n865), .ZN(n861) );
  OAI221_X1 U2836 ( .B1(n2103), .B2(n9489), .C1(n8406), .C2(n9486), .A(n883), 
        .ZN(n862) );
  NOR4_X1 U2837 ( .A1(n948), .A2(n949), .A3(n950), .A4(n951), .ZN(n947) );
  OAI221_X1 U2838 ( .B1(n2127), .B2(n9489), .C1(n8403), .C2(n9486), .A(n955), 
        .ZN(n948) );
  NOR4_X1 U2839 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1019)
         );
  OAI221_X1 U2840 ( .B1(n2159), .B2(n9489), .C1(n8399), .C2(n9486), .A(n1027), 
        .ZN(n1020) );
  NOR4_X1 U2841 ( .A1(n1398), .A2(n1399), .A3(n1400), .A4(n1401), .ZN(n1397)
         );
  OAI221_X1 U2842 ( .B1(n8474), .B2(n9511), .C1(n8238), .C2(n9508), .A(n1403), 
        .ZN(n1400) );
  NOR4_X1 U2843 ( .A1(n1200), .A2(n1201), .A3(n1202), .A4(n1203), .ZN(n1199)
         );
  OAI221_X1 U2844 ( .B1(n8253), .B2(n9512), .C1(n8216), .C2(n9509), .A(n1205), 
        .ZN(n1202) );
  NOR4_X1 U2845 ( .A1(n1272), .A2(n1273), .A3(n1274), .A4(n1275), .ZN(n1271)
         );
  OAI221_X1 U2846 ( .B1(n8249), .B2(n9511), .C1(n8224), .C2(n9508), .A(n1277), 
        .ZN(n1274) );
  NOR4_X1 U2847 ( .A1(n1128), .A2(n1129), .A3(n1130), .A4(n1131), .ZN(n1127)
         );
  OAI221_X1 U2848 ( .B1(n8257), .B2(n9512), .C1(n8208), .C2(n9509), .A(n1133), 
        .ZN(n1130) );
  NOR4_X1 U2849 ( .A1(n930), .A2(n931), .A3(n932), .A4(n933), .ZN(n929) );
  OAI221_X1 U2850 ( .B1(n2119), .B2(n9489), .C1(n8404), .C2(n9486), .A(n937), 
        .ZN(n930) );
  AND3_X1 U2851 ( .A1(ADD_RD2[1]), .A2(n10664), .A3(ADD_RD2[2]), .ZN(n2079) );
  AND3_X1 U2852 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[0]), .A3(ADD_RD2[2]), .ZN(n2078) );
  INV_X1 U2853 ( .A(ADD_WR[0]), .ZN(n9921) );
  INV_X1 U2854 ( .A(ADD_WR[2]), .ZN(n9919) );
  INV_X1 U2855 ( .A(ADD_WR[1]), .ZN(n9920) );
  NOR4_X1 U2856 ( .A1(n1344), .A2(n1345), .A3(n1346), .A4(n1347), .ZN(n1343)
         );
  OAI221_X1 U2857 ( .B1(n8924), .B2(n9439), .C1(n8892), .C2(n9436), .A(n1359), 
        .ZN(n1352) );
  AND3_X1 U2858 ( .A1(ADD_RD1[0]), .A2(n10659), .A3(ADD_RD1[2]), .ZN(n1467) );
  INV_X1 U2859 ( .A(ADD_RD2[1]), .ZN(n10663) );
  INV_X1 U2860 ( .A(ADD_RD2[0]), .ZN(n10664) );
  NOR4_X1 U2861 ( .A1(n1074), .A2(n1075), .A3(n1076), .A4(n1077), .ZN(n1073)
         );
  NOR4_X1 U2862 ( .A1(n1082), .A2(n1083), .A3(n1084), .A4(n1085), .ZN(n1072)
         );
  OAI221_X1 U2863 ( .B1(n8260), .B2(n9512), .C1(n8202), .C2(n9509), .A(n1079), 
        .ZN(n1076) );
  NOR4_X1 U2864 ( .A1(n1326), .A2(n1327), .A3(n1328), .A4(n1329), .ZN(n1325)
         );
  NOR4_X1 U2865 ( .A1(n1334), .A2(n1335), .A3(n1336), .A4(n1337), .ZN(n1324)
         );
  OAI221_X1 U2866 ( .B1(n8246), .B2(n9511), .C1(n8230), .C2(n9508), .A(n1331), 
        .ZN(n1328) );
  NOR4_X1 U2867 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1091)
         );
  NOR4_X1 U2868 ( .A1(n1100), .A2(n1101), .A3(n1102), .A4(n1103), .ZN(n1090)
         );
  OAI221_X1 U2869 ( .B1(n8259), .B2(n9512), .C1(n8204), .C2(n9509), .A(n1097), 
        .ZN(n1094) );
  AND3_X1 U2870 ( .A1(n10664), .A2(n10663), .A3(ADD_RD2[2]), .ZN(n2081) );
  AND3_X1 U2871 ( .A1(ADD_RD2[0]), .A2(n10663), .A3(ADD_RD2[2]), .ZN(n2080) );
  AND3_X1 U2872 ( .A1(n10660), .A2(n10659), .A3(ADD_RD1[2]), .ZN(n1466) );
  NAND2_X1 U2873 ( .A1(n1000), .A2(n1001), .ZN(N715) );
  NOR4_X1 U2874 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n1001)
         );
  NOR4_X1 U2875 ( .A1(n1010), .A2(n1011), .A3(n1012), .A4(n1013), .ZN(n1000)
         );
  OAI221_X1 U2876 ( .B1(n2151), .B2(n9489), .C1(n8400), .C2(n9486), .A(n1009), 
        .ZN(n1002) );
  NAND2_X1 U2877 ( .A1(n1378), .A2(n1379), .ZN(N694) );
  NOR4_X1 U2878 ( .A1(n1380), .A2(n1381), .A3(n1382), .A4(n1383), .ZN(n1379)
         );
  NOR4_X1 U2879 ( .A1(n1388), .A2(n1389), .A3(n1390), .A4(n1391), .ZN(n1378)
         );
  OAI221_X1 U2880 ( .B1(n8475), .B2(n9511), .C1(n8236), .C2(n9508), .A(n1385), 
        .ZN(n1382) );
  NAND2_X1 U2881 ( .A1(n1180), .A2(n1181), .ZN(N705) );
  NOR4_X1 U2882 ( .A1(n1182), .A2(n1183), .A3(n1184), .A4(n1185), .ZN(n1181)
         );
  NOR4_X1 U2883 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1180)
         );
  OAI221_X1 U2884 ( .B1(n8254), .B2(n9512), .C1(n8214), .C2(n9509), .A(n1187), 
        .ZN(n1184) );
  NAND2_X1 U2885 ( .A1(n1252), .A2(n1253), .ZN(N701) );
  NOR4_X1 U2886 ( .A1(n1254), .A2(n1255), .A3(n1256), .A4(n1257), .ZN(n1253)
         );
  NOR4_X1 U2887 ( .A1(n1262), .A2(n1263), .A3(n1264), .A4(n1265), .ZN(n1252)
         );
  OAI221_X1 U2888 ( .B1(n8250), .B2(n9511), .C1(n8222), .C2(n9508), .A(n1259), 
        .ZN(n1256) );
  NAND2_X1 U2889 ( .A1(n1108), .A2(n1109), .ZN(N709) );
  NOR4_X1 U2890 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .ZN(n1109)
         );
  NOR4_X1 U2891 ( .A1(n1118), .A2(n1119), .A3(n1120), .A4(n1121), .ZN(n1108)
         );
  OAI221_X1 U2892 ( .B1(n8258), .B2(n9512), .C1(n8206), .C2(n9509), .A(n1115), 
        .ZN(n1112) );
  NAND2_X1 U2893 ( .A1(n1414), .A2(n1415), .ZN(N692) );
  NOR4_X1 U2894 ( .A1(n1416), .A2(n1417), .A3(n1418), .A4(n1419), .ZN(n1415)
         );
  NOR4_X1 U2895 ( .A1(n1424), .A2(n1425), .A3(n1426), .A4(n1427), .ZN(n1414)
         );
  OAI221_X1 U2896 ( .B1(n8473), .B2(n9511), .C1(n8240), .C2(n9508), .A(n1421), 
        .ZN(n1418) );
  NAND2_X1 U2897 ( .A1(n1360), .A2(n1361), .ZN(N695) );
  NOR4_X1 U2898 ( .A1(n1362), .A2(n1363), .A3(n1364), .A4(n1365), .ZN(n1361)
         );
  NOR4_X1 U2899 ( .A1(n1370), .A2(n1371), .A3(n1372), .A4(n1373), .ZN(n1360)
         );
  OAI221_X1 U2900 ( .B1(n8476), .B2(n9511), .C1(n8234), .C2(n9508), .A(n1367), 
        .ZN(n1364) );
  NAND2_X1 U2901 ( .A1(n1162), .A2(n1163), .ZN(N706) );
  NOR4_X1 U2902 ( .A1(n1164), .A2(n1165), .A3(n1166), .A4(n1167), .ZN(n1163)
         );
  NOR4_X1 U2903 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1162)
         );
  OAI221_X1 U2904 ( .B1(n8255), .B2(n9512), .C1(n8212), .C2(n9509), .A(n1169), 
        .ZN(n1166) );
  NAND2_X1 U2905 ( .A1(n1234), .A2(n1235), .ZN(N702) );
  NOR4_X1 U2906 ( .A1(n1236), .A2(n1237), .A3(n1238), .A4(n1239), .ZN(n1235)
         );
  NOR4_X1 U2907 ( .A1(n1244), .A2(n1245), .A3(n1246), .A4(n1247), .ZN(n1234)
         );
  OAI221_X1 U2908 ( .B1(n8251), .B2(n9512), .C1(n8220), .C2(n9509), .A(n1241), 
        .ZN(n1238) );
  NAND2_X1 U2909 ( .A1(n1432), .A2(n1433), .ZN(N691) );
  NOR4_X1 U2910 ( .A1(n1434), .A2(n1435), .A3(n1436), .A4(n1437), .ZN(n1433)
         );
  NOR4_X1 U2911 ( .A1(n1442), .A2(n1443), .A3(n1444), .A4(n1445), .ZN(n1432)
         );
  OAI221_X1 U2912 ( .B1(n8472), .B2(n9511), .C1(n8242), .C2(n9508), .A(n1439), 
        .ZN(n1436) );
  NAND2_X1 U2913 ( .A1(n910), .A2(n911), .ZN(N720) );
  NOR4_X1 U2914 ( .A1(n912), .A2(n913), .A3(n914), .A4(n915), .ZN(n911) );
  NOR4_X1 U2915 ( .A1(n920), .A2(n921), .A3(n922), .A4(n923), .ZN(n910) );
  OAI221_X1 U2916 ( .B1(n2111), .B2(n9489), .C1(n8405), .C2(n9486), .A(n919), 
        .ZN(n912) );
  NAND2_X1 U2917 ( .A1(n964), .A2(n965), .ZN(N717) );
  NOR4_X1 U2918 ( .A1(n966), .A2(n967), .A3(n968), .A4(n969), .ZN(n965) );
  NOR4_X1 U2919 ( .A1(n974), .A2(n975), .A3(n976), .A4(n977), .ZN(n964) );
  OAI221_X1 U2920 ( .B1(n2135), .B2(n9489), .C1(n8402), .C2(n9486), .A(n973), 
        .ZN(n966) );
  NAND2_X1 U2921 ( .A1(n1036), .A2(n1037), .ZN(N713) );
  NOR4_X1 U2922 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1037)
         );
  NOR4_X1 U2923 ( .A1(n1046), .A2(n1047), .A3(n1048), .A4(n1049), .ZN(n1036)
         );
  OAI221_X1 U2924 ( .B1(n8262), .B2(n9512), .C1(n8198), .C2(n9509), .A(n1043), 
        .ZN(n1040) );
  NAND2_X1 U2925 ( .A1(n1288), .A2(n1289), .ZN(N699) );
  NOR4_X1 U2926 ( .A1(n1290), .A2(n1291), .A3(n1292), .A4(n1293), .ZN(n1289)
         );
  NOR4_X1 U2927 ( .A1(n1298), .A2(n1299), .A3(n1300), .A4(n1301), .ZN(n1288)
         );
  OAI221_X1 U2928 ( .B1(n8248), .B2(n9511), .C1(n8226), .C2(n9508), .A(n1295), 
        .ZN(n1292) );
  NAND2_X1 U2929 ( .A1(n1054), .A2(n1055), .ZN(N712) );
  NOR4_X1 U2930 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055)
         );
  NOR4_X1 U2931 ( .A1(n1064), .A2(n1065), .A3(n1066), .A4(n1067), .ZN(n1054)
         );
  OAI221_X1 U2932 ( .B1(n8261), .B2(n9512), .C1(n8200), .C2(n9509), .A(n1061), 
        .ZN(n1058) );
  AND3_X1 U2933 ( .A1(ENABLE), .A2(n9879), .A3(WR), .ZN(n849) );
  INV_X1 U2934 ( .A(ADD_RD1[0]), .ZN(n10660) );
  NAND2_X1 U2935 ( .A1(n2070), .A2(n2071), .ZN(N1020) );
  NOR4_X1 U2936 ( .A1(n2072), .A2(n2073), .A3(n2074), .A4(n2075), .ZN(n2071)
         );
  NAND2_X1 U2937 ( .A1(n2052), .A2(n2053), .ZN(N1021) );
  NOR4_X1 U2938 ( .A1(n2054), .A2(n2055), .A3(n2056), .A4(n2057), .ZN(n2053)
         );
  NAND2_X1 U2939 ( .A1(n2034), .A2(n2035), .ZN(N1022) );
  NOR4_X1 U2940 ( .A1(n2036), .A2(n2037), .A3(n2038), .A4(n2039), .ZN(n2035)
         );
  NAND2_X1 U2941 ( .A1(n2016), .A2(n2017), .ZN(N1023) );
  NOR4_X1 U2942 ( .A1(n2018), .A2(n2019), .A3(n2020), .A4(n2021), .ZN(n2017)
         );
  NAND2_X1 U2943 ( .A1(n1998), .A2(n1999), .ZN(N1024) );
  NOR4_X1 U2944 ( .A1(n2000), .A2(n2001), .A3(n2002), .A4(n2003), .ZN(n1999)
         );
  NAND2_X1 U2945 ( .A1(n1980), .A2(n1981), .ZN(N1025) );
  NOR4_X1 U2946 ( .A1(n1982), .A2(n1983), .A3(n1984), .A4(n1985), .ZN(n1981)
         );
  NAND2_X1 U2947 ( .A1(n1962), .A2(n1963), .ZN(N1026) );
  NOR4_X1 U2948 ( .A1(n1964), .A2(n1965), .A3(n1966), .A4(n1967), .ZN(n1963)
         );
  INV_X1 U2949 ( .A(DATAIN[3]), .ZN(n9913) );
  INV_X1 U2950 ( .A(DATAIN[4]), .ZN(n9912) );
  INV_X1 U2951 ( .A(DATAIN[5]), .ZN(n9911) );
  INV_X1 U2952 ( .A(DATAIN[6]), .ZN(n9910) );
  INV_X1 U2953 ( .A(DATAIN[7]), .ZN(n9909) );
  INV_X1 U2954 ( .A(DATAIN[8]), .ZN(n9908) );
  INV_X1 U2955 ( .A(DATAIN[31]), .ZN(n9885) );
  INV_X1 U2956 ( .A(DATAIN[0]), .ZN(n9916) );
  INV_X1 U2957 ( .A(DATAIN[1]), .ZN(n9915) );
  INV_X1 U2958 ( .A(DATAIN[2]), .ZN(n9914) );
  INV_X1 U2959 ( .A(DATAIN[10]), .ZN(n9906) );
  INV_X1 U2960 ( .A(DATAIN[11]), .ZN(n9905) );
  INV_X1 U2961 ( .A(DATAIN[12]), .ZN(n9904) );
  INV_X1 U2962 ( .A(DATAIN[13]), .ZN(n9903) );
  INV_X1 U2963 ( .A(DATAIN[14]), .ZN(n9902) );
  INV_X1 U2964 ( .A(DATAIN[15]), .ZN(n9901) );
  INV_X1 U2965 ( .A(DATAIN[16]), .ZN(n9900) );
  INV_X1 U2966 ( .A(DATAIN[17]), .ZN(n9899) );
  INV_X1 U2967 ( .A(DATAIN[18]), .ZN(n9898) );
  INV_X1 U2968 ( .A(DATAIN[19]), .ZN(n9897) );
  INV_X1 U2969 ( .A(DATAIN[20]), .ZN(n9896) );
  INV_X1 U2970 ( .A(DATAIN[21]), .ZN(n9895) );
  INV_X1 U2971 ( .A(DATAIN[22]), .ZN(n9894) );
  INV_X1 U2972 ( .A(DATAIN[23]), .ZN(n9893) );
  INV_X1 U2973 ( .A(DATAIN[24]), .ZN(n9892) );
  INV_X1 U2974 ( .A(DATAIN[25]), .ZN(n9891) );
  INV_X1 U2975 ( .A(DATAIN[26]), .ZN(n9890) );
  INV_X1 U2976 ( .A(DATAIN[27]), .ZN(n9889) );
  INV_X1 U2977 ( .A(DATAIN[28]), .ZN(n9888) );
  INV_X1 U2978 ( .A(DATAIN[29]), .ZN(n9887) );
  INV_X1 U2979 ( .A(DATAIN[30]), .ZN(n9886) );
  INV_X1 U2980 ( .A(DATAIN[9]), .ZN(n9907) );
  INV_X1 U2981 ( .A(ADD_RD2[3]), .ZN(n10662) );
  INV_X1 U2982 ( .A(ADD_RD2[4]), .ZN(n10661) );
  INV_X1 U2983 ( .A(ADD_RD1[3]), .ZN(n10658) );
  NAND2_X1 U2984 ( .A1(n1944), .A2(n1945), .ZN(N1027) );
  NOR4_X1 U2985 ( .A1(n1946), .A2(n1947), .A3(n1948), .A4(n1949), .ZN(n1945)
         );
  NAND2_X1 U2986 ( .A1(n1926), .A2(n1927), .ZN(N1028) );
  NOR4_X1 U2987 ( .A1(n1936), .A2(n1937), .A3(n1938), .A4(n1939), .ZN(n1926)
         );
  NAND2_X1 U2988 ( .A1(n1908), .A2(n1909), .ZN(N1029) );
  NOR4_X1 U2989 ( .A1(n1918), .A2(n1919), .A3(n1920), .A4(n1921), .ZN(n1908)
         );
  NAND2_X1 U2990 ( .A1(n1890), .A2(n1891), .ZN(N1030) );
  NOR4_X1 U2991 ( .A1(n1900), .A2(n1901), .A3(n1902), .A4(n1903), .ZN(n1890)
         );
  NAND2_X1 U2992 ( .A1(n1872), .A2(n1873), .ZN(N1031) );
  NOR4_X1 U2993 ( .A1(n1882), .A2(n1883), .A3(n1884), .A4(n1885), .ZN(n1872)
         );
  NAND2_X1 U2994 ( .A1(n1854), .A2(n1855), .ZN(N1032) );
  NOR4_X1 U2995 ( .A1(n1864), .A2(n1865), .A3(n1866), .A4(n1867), .ZN(n1854)
         );
  NAND2_X1 U2996 ( .A1(n1836), .A2(n1837), .ZN(N1033) );
  NOR4_X1 U2997 ( .A1(n1846), .A2(n1847), .A3(n1848), .A4(n1849), .ZN(n1836)
         );
  NAND2_X1 U2998 ( .A1(n1818), .A2(n1819), .ZN(N1034) );
  NOR4_X1 U2999 ( .A1(n1828), .A2(n1829), .A3(n1830), .A4(n1831), .ZN(n1818)
         );
  NAND2_X1 U3000 ( .A1(n1800), .A2(n1801), .ZN(N1035) );
  NOR4_X1 U3001 ( .A1(n1810), .A2(n1811), .A3(n1812), .A4(n1813), .ZN(n1800)
         );
  NAND2_X1 U3002 ( .A1(n1782), .A2(n1783), .ZN(N1036) );
  NOR4_X1 U3003 ( .A1(n1792), .A2(n1793), .A3(n1794), .A4(n1795), .ZN(n1782)
         );
  NAND2_X1 U3004 ( .A1(n1764), .A2(n1765), .ZN(N1037) );
  NOR4_X1 U3005 ( .A1(n1774), .A2(n1775), .A3(n1776), .A4(n1777), .ZN(n1764)
         );
  NAND2_X1 U3006 ( .A1(n1746), .A2(n1747), .ZN(N1038) );
  NOR4_X1 U3007 ( .A1(n1756), .A2(n1757), .A3(n1758), .A4(n1759), .ZN(n1746)
         );
  NAND2_X1 U3008 ( .A1(n1728), .A2(n1729), .ZN(N1039) );
  NOR4_X1 U3009 ( .A1(n1738), .A2(n1739), .A3(n1740), .A4(n1741), .ZN(n1728)
         );
  NAND2_X1 U3010 ( .A1(n1710), .A2(n1711), .ZN(N1040) );
  NOR4_X1 U3011 ( .A1(n1720), .A2(n1721), .A3(n1722), .A4(n1723), .ZN(n1710)
         );
  NAND2_X1 U3012 ( .A1(n1692), .A2(n1693), .ZN(N1041) );
  NOR4_X1 U3013 ( .A1(n1702), .A2(n1703), .A3(n1704), .A4(n1705), .ZN(n1692)
         );
  NAND2_X1 U3014 ( .A1(n1674), .A2(n1675), .ZN(N1042) );
  NOR4_X1 U3015 ( .A1(n1684), .A2(n1685), .A3(n1686), .A4(n1687), .ZN(n1674)
         );
  NAND2_X1 U3016 ( .A1(n1656), .A2(n1657), .ZN(N1043) );
  NOR4_X1 U3017 ( .A1(n1666), .A2(n1667), .A3(n1668), .A4(n1669), .ZN(n1656)
         );
  INV_X1 U3018 ( .A(ADD_WR[4]), .ZN(n9917) );
  INV_X1 U3019 ( .A(ADD_WR[3]), .ZN(n9918) );
  OAI221_X1 U3020 ( .B1(n8667), .B2(n9476), .C1(n8643), .C2(n9473), .A(n1230), 
        .ZN(n1229) );
  OAI221_X1 U3021 ( .B1(n8787), .B2(n9464), .C1(n8219), .C2(n9461), .A(n1231), 
        .ZN(n1228) );
  OAI221_X1 U3022 ( .B1(n8671), .B2(n9476), .C1(n8647), .C2(n9473), .A(n1158), 
        .ZN(n1157) );
  OAI221_X1 U3023 ( .B1(n8791), .B2(n9464), .C1(n8211), .C2(n9461), .A(n1159), 
        .ZN(n1156) );
  OAI221_X1 U3024 ( .B1(n8598), .B2(n9523), .C1(n8566), .C2(n9520), .A(n1456), 
        .ZN(n1455) );
  AOI22_X1 U3025 ( .A1(n9517), .A2(n10473), .B1(n9516), .B2(n10289), .ZN(n1456) );
  NAND2_X1 U3026 ( .A1(n1270), .A2(n1271), .ZN(N700) );
  NOR4_X1 U3027 ( .A1(n1280), .A2(n1281), .A3(n1282), .A4(n1283), .ZN(n1270)
         );
  NAND2_X1 U3028 ( .A1(n928), .A2(n929), .ZN(N719) );
  NOR4_X1 U3029 ( .A1(n938), .A2(n939), .A3(n940), .A4(n941), .ZN(n928) );
  NAND2_X1 U3030 ( .A1(n1324), .A2(n1325), .ZN(N697) );
  NAND2_X1 U3031 ( .A1(n1018), .A2(n1019), .ZN(N714) );
  NOR4_X1 U3032 ( .A1(n1028), .A2(n1029), .A3(n1030), .A4(n1031), .ZN(n1018)
         );
  NAND2_X1 U3033 ( .A1(n1090), .A2(n1091), .ZN(N710) );
  NAND2_X1 U3034 ( .A1(n1072), .A2(n1073), .ZN(N711) );
  OAI221_X1 U3035 ( .B1(n8654), .B2(n9475), .C1(n8630), .C2(n9472), .A(n1475), 
        .ZN(n1474) );
  OAI221_X1 U3036 ( .B1(n8774), .B2(n9463), .C1(n8245), .C2(n9460), .A(n1476), 
        .ZN(n1473) );
  NAND2_X1 U3037 ( .A1(n1198), .A2(n1199), .ZN(N704) );
  NOR4_X1 U3038 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1198)
         );
  NAND2_X1 U3039 ( .A1(n1126), .A2(n1127), .ZN(N708) );
  NOR4_X1 U3040 ( .A1(n1136), .A2(n1137), .A3(n1138), .A4(n1139), .ZN(n1126)
         );
  NAND2_X1 U3041 ( .A1(n946), .A2(n947), .ZN(N718) );
  NOR4_X1 U3042 ( .A1(n956), .A2(n957), .A3(n958), .A4(n959), .ZN(n946) );
  NAND2_X1 U3043 ( .A1(n860), .A2(n861), .ZN(N721) );
  NOR4_X1 U3044 ( .A1(n886), .A2(n887), .A3(n888), .A4(n889), .ZN(n860) );
  NAND2_X1 U3045 ( .A1(n1396), .A2(n1397), .ZN(N693) );
  NOR4_X1 U3046 ( .A1(n1406), .A2(n1407), .A3(n1408), .A4(n1409), .ZN(n1396)
         );
  NAND2_X1 U3047 ( .A1(n1216), .A2(n1217), .ZN(N703) );
  NOR4_X1 U3048 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1216)
         );
  NAND2_X1 U3049 ( .A1(n1144), .A2(n1145), .ZN(N707) );
  NOR4_X1 U3050 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1144)
         );
  NAND2_X1 U3051 ( .A1(n1450), .A2(n1451), .ZN(N690) );
  NOR4_X1 U3052 ( .A1(n1471), .A2(n1472), .A3(n1473), .A4(n1474), .ZN(n1450)
         );
  AND3_X1 U3053 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[0]), .A3(ADD_RD1[2]), .ZN(n1464) );
  AND3_X1 U3054 ( .A1(ADD_RD1[1]), .A2(n10660), .A3(ADD_RD1[2]), .ZN(n1468) );
  NOR3_X1 U3055 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(ADD_RD1[0]), .ZN(n1457) );
  NOR3_X1 U3056 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n10660), .ZN(n1459) );
  INV_X1 U3057 ( .A(ADD_RD1[1]), .ZN(n10659) );
  INV_X1 U3058 ( .A(ADD_RD1[4]), .ZN(n10665) );
  NOR4_X1 U3059 ( .A1(n1352), .A2(n1353), .A3(n1354), .A4(n1355), .ZN(n1342)
         );
  OAI221_X1 U3060 ( .B1(n8660), .B2(n9475), .C1(n8636), .C2(n9472), .A(n1356), 
        .ZN(n1355) );
  OAI221_X1 U3061 ( .B1(n8780), .B2(n9463), .C1(n8233), .C2(n9460), .A(n1357), 
        .ZN(n1354) );
  NAND2_X1 U3062 ( .A1(n1342), .A2(n1343), .ZN(N696) );
  NAND2_X1 U3063 ( .A1(n1306), .A2(n1307), .ZN(N698) );
  CLKBUF_X1 U3064 ( .A(n9882), .Z(n9877) );
  CLKBUF_X1 U3065 ( .A(n9881), .Z(n9878) );
  CLKBUF_X1 U3066 ( .A(n9880), .Z(n9879) );
endmodule


module DecodeUnit_DW01_add_0 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [9:1] carry;

  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XOR2_X1 U3 ( .A(A[6]), .B(B[6]), .Z(n3) );
  XOR2_X1 U4 ( .A(n3), .B(carry[6]), .Z(SUM[6]) );
  NAND3_X1 U8 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[7]) );
  XOR2_X1 U9 ( .A(A[7]), .B(B[7]), .Z(n7) );
  XOR2_X1 U10 ( .A(n7), .B(carry[7]), .Z(SUM[7]) );
  NAND3_X1 U14 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[8]) );
  XOR2_X1 U15 ( .A(B[1]), .B(A[1]), .Z(n11) );
  XOR2_X1 U16 ( .A(n2), .B(n11), .Z(SUM[1]) );
  NAND3_X1 U20 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[2]) );
  XOR2_X1 U21 ( .A(B[2]), .B(A[2]), .Z(n15) );
  XOR2_X1 U22 ( .A(carry[2]), .B(n15), .Z(SUM[2]) );
  NAND3_X1 U26 ( .A1(n16), .A2(n17), .A3(n18), .ZN(carry[3]) );
  XOR2_X1 U27 ( .A(B[9]), .B(A[9]), .Z(n19) );
  XOR2_X1 U28 ( .A(carry[9]), .B(n19), .Z(SUM[9]) );
  NAND2_X1 U2 ( .A1(B[7]), .A2(carry[7]), .ZN(n10) );
  NAND2_X1 U5 ( .A1(A[6]), .A2(B[6]), .ZN(n4) );
  NAND2_X1 U6 ( .A1(A[6]), .A2(carry[6]), .ZN(n5) );
  NAND2_X1 U7 ( .A1(B[6]), .A2(carry[6]), .ZN(n6) );
  NAND2_X1 U11 ( .A1(B[1]), .A2(A[1]), .ZN(n14) );
  NAND2_X1 U12 ( .A1(n2), .A2(B[1]), .ZN(n12) );
  NAND2_X1 U13 ( .A1(n2), .A2(A[1]), .ZN(n13) );
  NAND2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n18) );
  NAND2_X1 U18 ( .A1(carry[2]), .A2(B[2]), .ZN(n16) );
  AND2_X1 U19 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
  NAND2_X1 U23 ( .A1(A[7]), .A2(B[7]), .ZN(n8) );
  NAND2_X1 U24 ( .A1(A[7]), .A2(carry[7]), .ZN(n9) );
  NAND2_X1 U25 ( .A1(carry[2]), .A2(A[2]), .ZN(n17) );
endmodule


module DecodeUnit ( clock, reset, JMP, RegDestination, en2, SignSelect, 
        BranchCondSel, BRANCHenable, RD1, RD2, WR, Instruction, ADD_WR, DATAIN, 
        NPCfromIF, OUT1, OUT2, OUTNPC, OUTIMM, NPCtoEX, AddressWtoEX, 
        BRANCHtoFetch );
  input [31:0] Instruction;
  input [4:0] ADD_WR;
  input [31:0] DATAIN;
  input [31:0] NPCfromIF;
  output [31:0] OUT1;
  output [31:0] OUT2;
  output [31:0] OUTNPC;
  output [31:0] OUTIMM;
  output [31:0] NPCtoEX;
  output [31:0] AddressWtoEX;
  input clock, reset, JMP, RegDestination, en2, SignSelect, BranchCondSel,
         BRANCHenable, RD1, RD2, WR;
  output BRANCHtoFetch;
  wire   BranchTaken, n4, n20;
  wire   [31:0] AddressW;
  wire   [31:0] MuxtoIMM;
  wire   [31:0] RFOUT1;
  wire   [31:0] RFOUT2;
  assign OUTNPC[10] = 1'b0;
  assign OUTNPC[11] = 1'b0;
  assign OUTNPC[12] = 1'b0;
  assign OUTNPC[13] = 1'b0;
  assign OUTNPC[14] = 1'b0;
  assign OUTNPC[15] = 1'b0;
  assign OUTNPC[16] = 1'b0;
  assign OUTNPC[17] = 1'b0;
  assign OUTNPC[18] = 1'b0;
  assign OUTNPC[19] = 1'b0;
  assign OUTNPC[20] = 1'b0;
  assign OUTNPC[21] = 1'b0;
  assign OUTNPC[22] = 1'b0;
  assign OUTNPC[23] = 1'b0;
  assign OUTNPC[24] = 1'b0;
  assign OUTNPC[25] = 1'b0;
  assign OUTNPC[26] = 1'b0;
  assign OUTNPC[27] = 1'b0;
  assign OUTNPC[28] = 1'b0;
  assign OUTNPC[29] = 1'b0;
  assign OUTNPC[30] = 1'b0;
  assign OUTNPC[31] = 1'b0;

  Mux41 ADDRESS_MUX ( .a({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Instruction[20:16]}), .b({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, Instruction[15:11]}), .c({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1}), .d({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .sel({JMP, RegDestination}), .y(AddressW) );
  Mux21_5 MUX ( .a({Instruction[15], Instruction[15], Instruction[15], 
        Instruction[15], Instruction[15], Instruction[15], Instruction[15], 
        Instruction[15], Instruction[15], Instruction[15], Instruction[15], 
        Instruction[15], Instruction[15], Instruction[15], Instruction[15], 
        Instruction[15], Instruction[15:0]}), .b({n20, n20, n20, n20, n20, n20, 
        n20, Instruction[24:0]}), .sel(SignSelect), .y(MuxtoIMM) );
  BranchUnit BRANCH ( .a(RFOUT1), .sel(BranchCondSel), .y(BranchTaken) );
  reg_11 IMM_REG ( .clock(clock), .reset(reset), .load(en2), .i(MuxtoIMM), .o(
        OUTIMM) );
  reg_10 OUT1_REG ( .clock(clock), .reset(reset), .load(en2), .i(RFOUT1), .o(
        OUT1) );
  reg_9 OUT2_REG ( .clock(clock), .reset(reset), .load(en2), .i(RFOUT2), .o(
        OUT2) );
  reg_8 NXPC_REG ( .clock(clock), .reset(reset), .load(en2), .i(NPCfromIF), 
        .o(NPCtoEX) );
  reg_7 ADD_WR_REG ( .clock(clock), .reset(reset), .load(en2), .i(AddressW), 
        .o(AddressWtoEX) );
  register_file RF ( .CLK(clock), .RESET(reset), .ENABLE(1'b1), .RD1(RD1), 
        .RD2(RD2), .WR(WR), .ADD_WR(ADD_WR), .ADD_RD1(Instruction[25:21]), 
        .ADD_RD2(Instruction[20:16]), .DATAIN(DATAIN), .OUT1(RFOUT1), .OUT2(
        RFOUT2) );
  DecodeUnit_DW01_add_0 add_142 ( .A(NPCfromIF[9:0]), .B(MuxtoIMM[11:2]), .CI(
        1'b0), .SUM(OUTNPC[9:0]) );
  INV_X1 U3 ( .A(n4), .ZN(BRANCHtoFetch) );
  CLKBUF_X1 U5 ( .A(Instruction[25]), .Z(n20) );
  AOI21_X1 U6 ( .B1(BranchTaken), .B2(BRANCHenable), .A(JMP), .ZN(n4) );
endmodule


module Mux21_4 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, net131825, net131826, net131827, net131845, net133025,
         net133017, net133015, net133013, net133009, net133005, net133003,
         net133001, net141441, net141472, net141479, net141488, net141492,
         net141590, n42, n172, n173, n174, n175, n177, n178;
  assign y[10] = net131825;
  assign y[11] = net131826;
  assign y[12] = net131827;
  assign y[30] = net131845;

  CLKBUF_X1 U1 ( .A(net133009), .Z(net141590) );
  CLKBUF_X1 U2 ( .A(net141441), .Z(n172) );
  AOI22_X1 U3 ( .A1(net141479), .A2(a[30]), .B1(net133009), .B2(b[30]), .ZN(
        n42) );
  INV_X1 U4 ( .A(n42), .ZN(net131845) );
  BUF_X1 U5 ( .A(n174), .Z(n173) );
  AOI22_X1 U6 ( .A1(net133003), .A2(a[12]), .B1(n173), .B2(b[12]), .ZN(n62) );
  AOI22_X1 U7 ( .A1(net141492), .A2(a[11]), .B1(n173), .B2(b[11]), .ZN(n63) );
  AOI22_X1 U8 ( .A1(net133001), .A2(a[10]), .B1(net133017), .B2(b[10]), .ZN(
        n64) );
  INV_X1 U9 ( .A(sel), .ZN(n174) );
  BUF_X1 U10 ( .A(n174), .Z(net133005) );
  INV_X1 U11 ( .A(n174), .ZN(net133003) );
  INV_X1 U12 ( .A(n174), .ZN(net141492) );
  INV_X1 U13 ( .A(n175), .ZN(net141479) );
  INV_X1 U14 ( .A(sel), .ZN(n175) );
  BUF_X2 U15 ( .A(n175), .Z(net133009) );
  BUF_X2 U16 ( .A(n175), .Z(net133017) );
  INV_X1 U17 ( .A(sel), .ZN(net133025) );
  CLKBUF_X1 U18 ( .A(net141441), .Z(net141488) );
  BUF_X1 U19 ( .A(net133025), .Z(net133015) );
  INV_X1 U20 ( .A(net133025), .ZN(net133001) );
  INV_X1 U21 ( .A(net133003), .ZN(net141472) );
  INV_X1 U22 ( .A(net133025), .ZN(net141441) );
  OR2_X1 U23 ( .A1(n177), .A2(n178), .ZN(y[28]) );
  AND2_X1 U24 ( .A1(net133001), .A2(a[28]), .ZN(n177) );
  AND2_X1 U25 ( .A1(net133009), .A2(b[28]), .ZN(n178) );
  BUF_X1 U26 ( .A(net133025), .Z(net133013) );
  INV_X1 U27 ( .A(n43), .ZN(y[2]) );
  INV_X1 U28 ( .A(n54), .ZN(y[1]) );
  INV_X1 U29 ( .A(n40), .ZN(y[3]) );
  INV_X1 U30 ( .A(n39), .ZN(y[4]) );
  INV_X1 U31 ( .A(n38), .ZN(y[5]) );
  AOI22_X1 U32 ( .A1(a[4]), .A2(net141488), .B1(b[4]), .B2(net141472), .ZN(n39) );
  AOI22_X1 U33 ( .A1(a[5]), .A2(net141441), .B1(b[5]), .B2(net141590), .ZN(n38) );
  AOI22_X1 U34 ( .A1(a[3]), .A2(n172), .B1(b[3]), .B2(net141472), .ZN(n40) );
  AOI22_X1 U35 ( .A1(net141479), .A2(a[9]), .B1(n173), .B2(b[9]), .ZN(n34) );
  INV_X1 U36 ( .A(n36), .ZN(y[7]) );
  AOI22_X1 U37 ( .A1(a[7]), .A2(net133003), .B1(b[7]), .B2(net133013), .ZN(n36) );
  INV_X1 U38 ( .A(n34), .ZN(y[9]) );
  AOI22_X1 U39 ( .A1(a[6]), .A2(net141441), .B1(net133005), .B2(b[6]), .ZN(n37) );
  INV_X1 U40 ( .A(n57), .ZN(y[17]) );
  INV_X1 U41 ( .A(n46), .ZN(y[27]) );
  INV_X1 U42 ( .A(n52), .ZN(y[21]) );
  INV_X1 U43 ( .A(n56), .ZN(y[18]) );
  INV_X1 U44 ( .A(n47), .ZN(y[26]) );
  INV_X1 U45 ( .A(n55), .ZN(y[19]) );
  INV_X1 U46 ( .A(n59), .ZN(y[15]) );
  INV_X1 U47 ( .A(n44), .ZN(y[29]) );
  INV_X1 U48 ( .A(n65), .ZN(y[0]) );
  INV_X1 U49 ( .A(n35), .ZN(y[8]) );
  AOI22_X1 U50 ( .A1(a[8]), .A2(net133003), .B1(b[8]), .B2(net133005), .ZN(n35) );
  INV_X1 U51 ( .A(n58), .ZN(y[16]) );
  INV_X1 U52 ( .A(n53), .ZN(y[20]) );
  INV_X1 U53 ( .A(n63), .ZN(net131826) );
  INV_X1 U54 ( .A(n37), .ZN(y[6]) );
  INV_X1 U55 ( .A(n60), .ZN(y[14]) );
  INV_X1 U56 ( .A(n41), .ZN(y[31]) );
  INV_X1 U57 ( .A(n48), .ZN(y[25]) );
  INV_X1 U58 ( .A(n62), .ZN(net131827) );
  INV_X1 U59 ( .A(n49), .ZN(y[24]) );
  INV_X1 U60 ( .A(n50), .ZN(y[23]) );
  AOI22_X1 U61 ( .A1(a[31]), .A2(net141441), .B1(net133005), .B2(b[31]), .ZN(
        n41) );
  INV_X1 U62 ( .A(n61), .ZN(y[13]) );
  AOI22_X1 U63 ( .A1(a[2]), .A2(net141488), .B1(b[2]), .B2(net141472), .ZN(n43) );
  INV_X1 U64 ( .A(n51), .ZN(y[22]) );
  AOI22_X1 U65 ( .A1(net133003), .A2(a[27]), .B1(net133013), .B2(b[27]), .ZN(
        n46) );
  AOI22_X1 U66 ( .A1(a[26]), .A2(net141479), .B1(b[26]), .B2(net133017), .ZN(
        n47) );
  AOI22_X1 U67 ( .A1(net133001), .A2(a[29]), .B1(net133015), .B2(b[29]), .ZN(
        n44) );
  AOI22_X1 U68 ( .A1(a[20]), .A2(net133003), .B1(b[20]), .B2(net133017), .ZN(
        n53) );
  AOI22_X1 U69 ( .A1(net141479), .A2(a[21]), .B1(net133013), .B2(b[21]), .ZN(
        n52) );
  AOI22_X1 U70 ( .A1(net141479), .A2(a[25]), .B1(net133009), .B2(b[25]), .ZN(
        n48) );
  AOI22_X1 U71 ( .A1(net133001), .A2(a[24]), .B1(net133009), .B2(b[24]), .ZN(
        n49) );
  AOI22_X1 U72 ( .A1(net141479), .A2(a[23]), .B1(net133009), .B2(b[23]), .ZN(
        n50) );
  AOI22_X1 U73 ( .A1(net133001), .A2(a[22]), .B1(net133015), .B2(b[22]), .ZN(
        n51) );
  AOI22_X1 U74 ( .A1(a[1]), .A2(net141441), .B1(net141590), .B2(b[1]), .ZN(n54) );
  AOI22_X1 U75 ( .A1(a[0]), .A2(net141441), .B1(b[0]), .B2(net133017), .ZN(n65) );
  INV_X1 U76 ( .A(n64), .ZN(net131825) );
  AOI22_X1 U77 ( .A1(net141492), .A2(a[19]), .B1(n173), .B2(b[19]), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(net141492), .A2(a[18]), .B1(net133015), .B2(b[18]), .ZN(
        n56) );
  AOI22_X1 U79 ( .A1(a[17]), .A2(net141492), .B1(net133013), .B2(b[17]), .ZN(
        n57) );
  AOI22_X1 U80 ( .A1(a[14]), .A2(net133003), .B1(b[14]), .B2(net133017), .ZN(
        n60) );
  AOI22_X1 U81 ( .A1(net141492), .A2(a[16]), .B1(net133005), .B2(b[16]), .ZN(
        n58) );
  AOI22_X1 U82 ( .A1(net141441), .A2(a[15]), .B1(net133005), .B2(b[15]), .ZN(
        n59) );
  AOI22_X1 U83 ( .A1(net141492), .A2(a[13]), .B1(b[13]), .B2(net133017), .ZN(
        n61) );
endmodule


module Mux21_3 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249;

  INV_X1 U1 ( .A(n221), .ZN(y[12]) );
  INV_X1 U2 ( .A(n231), .ZN(y[21]) );
  INV_X1 U3 ( .A(n234), .ZN(y[24]) );
  INV_X1 U4 ( .A(n245), .ZN(y[5]) );
  INV_X1 U5 ( .A(n238), .ZN(y[28]) );
  INV_X1 U6 ( .A(n230), .ZN(y[20]) );
  INV_X1 U7 ( .A(n249), .ZN(y[9]) );
  INV_X1 U8 ( .A(n229), .ZN(y[1]) );
  INV_X1 U9 ( .A(n222), .ZN(y[13]) );
  INV_X1 U10 ( .A(n235), .ZN(y[25]) );
  INV_X1 U11 ( .A(n223), .ZN(y[14]) );
  INV_X1 U12 ( .A(n225), .ZN(y[16]) );
  INV_X1 U13 ( .A(n226), .ZN(y[17]) );
  INV_X1 U14 ( .A(n227), .ZN(y[18]) );
  INV_X1 U15 ( .A(n232), .ZN(y[22]) );
  INV_X1 U16 ( .A(n236), .ZN(y[26]) );
  INV_X1 U17 ( .A(n243), .ZN(y[3]) );
  INV_X1 U18 ( .A(n247), .ZN(y[7]) );
  INV_X1 U19 ( .A(n220), .ZN(y[11]) );
  INV_X1 U20 ( .A(n224), .ZN(y[15]) );
  INV_X1 U21 ( .A(n228), .ZN(y[19]) );
  INV_X1 U22 ( .A(n233), .ZN(y[23]) );
  INV_X1 U23 ( .A(n237), .ZN(y[27]) );
  INV_X2 U24 ( .A(n184), .ZN(n173) );
  MUX2_X1 U25 ( .A(b[0]), .B(a[0]), .S(sel), .Z(y[0]) );
  CLKBUF_X1 U26 ( .A(n185), .Z(n183) );
  CLKBUF_X1 U27 ( .A(n185), .Z(n182) );
  CLKBUF_X1 U28 ( .A(sel), .Z(n172) );
  INV_X1 U29 ( .A(n184), .ZN(n174) );
  BUF_X1 U30 ( .A(n186), .Z(n179) );
  BUF_X1 U31 ( .A(n186), .Z(n178) );
  BUF_X1 U32 ( .A(n186), .Z(n180) );
  BUF_X1 U33 ( .A(n186), .Z(n181) );
  BUF_X1 U34 ( .A(n185), .Z(n184) );
  BUF_X1 U35 ( .A(n186), .Z(n177) );
  BUF_X1 U36 ( .A(n186), .Z(n176) );
  INV_X1 U37 ( .A(n172), .ZN(n185) );
  INV_X1 U38 ( .A(n172), .ZN(n186) );
  INV_X1 U39 ( .A(n241), .ZN(y[30]) );
  AOI22_X1 U40 ( .A1(a[30]), .A2(n174), .B1(b[30]), .B2(n178), .ZN(n241) );
  AOI22_X1 U41 ( .A1(a[25]), .A2(n174), .B1(b[25]), .B2(n179), .ZN(n235) );
  AOI22_X1 U42 ( .A1(a[1]), .A2(n173), .B1(b[1]), .B2(n181), .ZN(n229) );
  AOI22_X1 U43 ( .A1(a[26]), .A2(n174), .B1(b[26]), .B2(n179), .ZN(n236) );
  AOI22_X1 U44 ( .A1(a[22]), .A2(n174), .B1(b[22]), .B2(n180), .ZN(n232) );
  AOI22_X1 U45 ( .A1(a[23]), .A2(n174), .B1(b[23]), .B2(n180), .ZN(n233) );
  INV_X1 U46 ( .A(n242), .ZN(y[31]) );
  AOI22_X1 U47 ( .A1(a[13]), .A2(n173), .B1(b[13]), .B2(n182), .ZN(n222) );
  AOI22_X1 U48 ( .A1(a[28]), .A2(n174), .B1(b[28]), .B2(n178), .ZN(n238) );
  AOI22_X1 U49 ( .A1(a[18]), .A2(n173), .B1(b[18]), .B2(n181), .ZN(n227) );
  AOI22_X1 U50 ( .A1(a[15]), .A2(n173), .B1(b[15]), .B2(n182), .ZN(n224) );
  AOI22_X1 U51 ( .A1(a[19]), .A2(n173), .B1(b[19]), .B2(n181), .ZN(n228) );
  AOI22_X1 U52 ( .A1(a[17]), .A2(n173), .B1(b[17]), .B2(n181), .ZN(n226) );
  AOI22_X1 U53 ( .A1(a[24]), .A2(n174), .B1(b[24]), .B2(n179), .ZN(n234) );
  AOI22_X1 U54 ( .A1(a[27]), .A2(n174), .B1(b[27]), .B2(n179), .ZN(n237) );
  AOI22_X1 U55 ( .A1(a[14]), .A2(n173), .B1(b[14]), .B2(n182), .ZN(n223) );
  AOI22_X1 U56 ( .A1(a[12]), .A2(n173), .B1(b[12]), .B2(n183), .ZN(n221) );
  AOI22_X1 U57 ( .A1(a[11]), .A2(n173), .B1(b[11]), .B2(n183), .ZN(n220) );
  AOI22_X1 U58 ( .A1(a[16]), .A2(n173), .B1(b[16]), .B2(n182), .ZN(n225) );
  AOI22_X1 U59 ( .A1(a[2]), .A2(n174), .B1(b[2]), .B2(n178), .ZN(n240) );
  INV_X1 U60 ( .A(n239), .ZN(y[29]) );
  AOI22_X1 U61 ( .A1(a[29]), .A2(n174), .B1(b[29]), .B2(n178), .ZN(n239) );
  AOI22_X1 U62 ( .A1(a[21]), .A2(n174), .B1(b[21]), .B2(n180), .ZN(n231) );
  AOI22_X1 U63 ( .A1(a[20]), .A2(n174), .B1(b[20]), .B2(n180), .ZN(n230) );
  AOI22_X1 U64 ( .A1(a[10]), .A2(n173), .B1(b[10]), .B2(n183), .ZN(n219) );
  AOI22_X1 U65 ( .A1(a[31]), .A2(n175), .B1(b[31]), .B2(n177), .ZN(n242) );
  AOI22_X1 U66 ( .A1(a[5]), .A2(n175), .B1(b[5]), .B2(n177), .ZN(n245) );
  AOI22_X1 U67 ( .A1(n175), .A2(a[9]), .B1(b[9]), .B2(n176), .ZN(n249) );
  AOI22_X1 U68 ( .A1(a[3]), .A2(n175), .B1(b[3]), .B2(n177), .ZN(n243) );
  AOI22_X1 U69 ( .A1(a[7]), .A2(n175), .B1(b[7]), .B2(n176), .ZN(n247) );
  AOI22_X1 U70 ( .A1(a[8]), .A2(n175), .B1(b[8]), .B2(n176), .ZN(n248) );
  AOI22_X1 U71 ( .A1(a[6]), .A2(n175), .B1(b[6]), .B2(n176), .ZN(n246) );
  AOI22_X1 U72 ( .A1(a[4]), .A2(n175), .B1(b[4]), .B2(n177), .ZN(n244) );
  INV_X1 U73 ( .A(n184), .ZN(n175) );
  INV_X2 U74 ( .A(n219), .ZN(y[10]) );
  INV_X2 U75 ( .A(n248), .ZN(y[8]) );
  INV_X2 U76 ( .A(n246), .ZN(y[6]) );
  INV_X2 U77 ( .A(n244), .ZN(y[4]) );
  INV_X2 U78 ( .A(n240), .ZN(y[2]) );
endmodule


module Mux21_2 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n43, n44, n45, net132218, net132244, net132245, net132246, net132961,
         net132955, net132953, net132951, net132949, net132947, net132943,
         net132941, net132937, net132935, n172, n173, n174, n175, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227;
  assign y[2] = net132218;
  assign y[28] = net132244;
  assign y[29] = net132245;
  assign y[30] = net132246;

  INV_X1 U1 ( .A(n174), .ZN(net132937) );
  INV_X1 U2 ( .A(n174), .ZN(net132935) );
  INV_X1 U3 ( .A(n213), .ZN(y[1]) );
  BUF_X1 U4 ( .A(n175), .Z(n174) );
  MUX2_X1 U5 ( .A(b[12]), .B(a[12]), .S(sel), .Z(y[12]) );
  MUX2_X1 U6 ( .A(b[16]), .B(a[16]), .S(sel), .Z(y[16]) );
  MUX2_X1 U7 ( .A(b[6]), .B(a[6]), .S(sel), .Z(y[6]) );
  MUX2_X1 U8 ( .A(b[24]), .B(a[24]), .S(sel), .Z(y[24]) );
  INV_X1 U9 ( .A(n43), .ZN(net132218) );
  AOI22_X1 U10 ( .A1(a[30]), .A2(net132937), .B1(b[30]), .B2(n173), .ZN(n172)
         );
  INV_X1 U11 ( .A(n172), .ZN(net132246) );
  BUF_X1 U12 ( .A(n175), .Z(n173) );
  AOI22_X1 U13 ( .A1(a[28]), .A2(net132937), .B1(b[28]), .B2(n173), .ZN(n45)
         );
  AOI22_X1 U14 ( .A1(a[2]), .A2(net132937), .B1(b[2]), .B2(n173), .ZN(n43) );
  AOI22_X1 U15 ( .A1(a[29]), .A2(net132937), .B1(b[29]), .B2(n173), .ZN(n44)
         );
  CLKBUF_X1 U16 ( .A(n175), .Z(net132943) );
  BUF_X1 U17 ( .A(net132961), .Z(net132941) );
  INV_X1 U18 ( .A(sel), .ZN(net132961) );
  INV_X1 U19 ( .A(sel), .ZN(n175) );
  BUF_X1 U20 ( .A(n175), .Z(net132953) );
  BUF_X1 U21 ( .A(n175), .Z(net132955) );
  INV_X1 U22 ( .A(n220), .ZN(y[27]) );
  INV_X1 U23 ( .A(n226), .ZN(y[8]) );
  INV_X1 U24 ( .A(n214), .ZN(y[20]) );
  INV_X1 U25 ( .A(n206), .ZN(y[11]) );
  INV_X1 U26 ( .A(n225), .ZN(y[7]) );
  INV_X1 U27 ( .A(n227), .ZN(y[9]) );
  INV_X1 U28 ( .A(n208), .ZN(y[14]) );
  INV_X1 U29 ( .A(n215), .ZN(y[21]) );
  INV_X1 U30 ( .A(n44), .ZN(net132245) );
  INV_X1 U31 ( .A(n209), .ZN(y[15]) );
  INV_X1 U32 ( .A(n45), .ZN(net132244) );
  INV_X1 U33 ( .A(n218), .ZN(y[25]) );
  INV_X1 U34 ( .A(n207), .ZN(y[13]) );
  INV_X1 U35 ( .A(n217), .ZN(y[23]) );
  INV_X1 U36 ( .A(n205), .ZN(y[10]) );
  INV_X1 U37 ( .A(n211), .ZN(y[18]) );
  INV_X1 U38 ( .A(n210), .ZN(y[17]) );
  BUF_X1 U39 ( .A(net132961), .Z(net132949) );
  BUF_X1 U40 ( .A(net132961), .Z(net132951) );
  BUF_X1 U41 ( .A(net132961), .Z(net132947) );
  AOI22_X1 U42 ( .A1(net132935), .A2(a[9]), .B1(b[9]), .B2(net132941), .ZN(
        n227) );
  INV_X1 U43 ( .A(n219), .ZN(y[26]) );
  AOI22_X1 U44 ( .A1(a[14]), .A2(net132935), .B1(b[14]), .B2(net132953), .ZN(
        n208) );
  AOI22_X1 U45 ( .A1(a[15]), .A2(net132935), .B1(b[15]), .B2(net132953), .ZN(
        n209) );
  INV_X1 U46 ( .A(n204), .ZN(y[0]) );
  AOI22_X1 U47 ( .A1(a[0]), .A2(net132935), .B1(b[0]), .B2(net132955), .ZN(
        n204) );
  AOI22_X1 U48 ( .A1(a[21]), .A2(net132937), .B1(b[21]), .B2(net132949), .ZN(
        n215) );
  AOI22_X1 U49 ( .A1(a[20]), .A2(net132937), .B1(b[20]), .B2(net132949), .ZN(
        n214) );
  AOI22_X1 U50 ( .A1(a[1]), .A2(net132935), .B1(b[1]), .B2(net132951), .ZN(
        n213) );
  INV_X1 U51 ( .A(n222), .ZN(y[3]) );
  AOI22_X1 U52 ( .A1(a[3]), .A2(net132937), .B1(b[3]), .B2(net132943), .ZN(
        n222) );
  INV_X1 U53 ( .A(n223), .ZN(y[4]) );
  AOI22_X1 U54 ( .A1(a[4]), .A2(net132935), .B1(b[4]), .B2(net132943), .ZN(
        n223) );
  INV_X1 U55 ( .A(n224), .ZN(y[5]) );
  AOI22_X1 U56 ( .A1(a[5]), .A2(net132937), .B1(b[5]), .B2(net132943), .ZN(
        n224) );
  AOI22_X1 U57 ( .A1(a[11]), .A2(net132935), .B1(b[11]), .B2(net132955), .ZN(
        n206) );
  INV_X1 U58 ( .A(n221), .ZN(y[31]) );
  INV_X1 U59 ( .A(n212), .ZN(y[19]) );
  AOI22_X1 U60 ( .A1(a[10]), .A2(net132935), .B1(b[10]), .B2(net132955), .ZN(
        n205) );
  AOI22_X1 U61 ( .A1(a[27]), .A2(net132937), .B1(b[27]), .B2(net132947), .ZN(
        n220) );
  AOI22_X1 U62 ( .A1(a[7]), .A2(net132935), .B1(b[7]), .B2(net132941), .ZN(
        n225) );
  INV_X1 U63 ( .A(n216), .ZN(y[22]) );
  AOI22_X1 U64 ( .A1(a[22]), .A2(net132937), .B1(b[22]), .B2(net132949), .ZN(
        n216) );
  AOI22_X1 U65 ( .A1(a[17]), .A2(net132935), .B1(b[17]), .B2(net132951), .ZN(
        n210) );
  AOI22_X1 U66 ( .A1(a[25]), .A2(net132937), .B1(b[25]), .B2(net132947), .ZN(
        n218) );
  AOI22_X1 U67 ( .A1(a[18]), .A2(net132935), .B1(b[18]), .B2(net132951), .ZN(
        n211) );
  AOI22_X1 U68 ( .A1(a[26]), .A2(net132937), .B1(b[26]), .B2(net132947), .ZN(
        n219) );
  AOI22_X1 U69 ( .A1(a[19]), .A2(net132935), .B1(b[19]), .B2(net132951), .ZN(
        n212) );
  AOI22_X1 U70 ( .A1(a[8]), .A2(net132937), .B1(b[8]), .B2(net132941), .ZN(
        n226) );
  AOI22_X1 U71 ( .A1(a[31]), .A2(net132935), .B1(b[31]), .B2(net132943), .ZN(
        n221) );
  AOI22_X1 U72 ( .A1(a[23]), .A2(net132937), .B1(b[23]), .B2(net132949), .ZN(
        n217) );
  AOI22_X1 U73 ( .A1(a[13]), .A2(net132935), .B1(b[13]), .B2(net132953), .ZN(
        n207) );
endmodule


module SHIFTER_M32_N5_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \temp_int_SH[4] , \SHMAG[5] , \MR_int[1][31] , \MR_int[1][30] ,
         \MR_int[1][29] , \MR_int[1][28] , \MR_int[1][27] , \MR_int[1][26] ,
         \MR_int[1][25] , \MR_int[1][24] , \MR_int[1][22] , \MR_int[1][21] ,
         \MR_int[1][16] , \MR_int[1][15] , \MR_int[1][14] , \MR_int[1][13] ,
         \MR_int[1][12] , \MR_int[1][11] , \MR_int[1][10] , \MR_int[1][9] ,
         \MR_int[1][8] , \MR_int[1][7] , \MR_int[1][6] , \MR_int[1][5] ,
         \MR_int[1][4] , \MR_int[1][3] , \MR_int[1][2] , \MR_int[1][1] ,
         \MR_int[2][31] , \MR_int[2][30] , \MR_int[2][29] , \MR_int[2][27] ,
         \MR_int[2][26] , \MR_int[2][25] , \MR_int[2][24] , \MR_int[2][23] ,
         \MR_int[2][22] , \MR_int[2][21] , \MR_int[2][20] , \MR_int[2][19] ,
         \MR_int[2][16] , \MR_int[2][15] , \MR_int[2][11] , \MR_int[2][10] ,
         \MR_int[2][9] , \MR_int[2][8] , \MR_int[2][7] , \MR_int[2][6] ,
         \MR_int[2][5] , \MR_int[2][4] , \MR_int[2][3] , \MR_int[2][2] ,
         \MR_int[2][1] , \MR_int[3][31] , \MR_int[3][30] , \MR_int[3][29] ,
         \MR_int[3][27] , \MR_int[3][26] , \MR_int[3][25] , \MR_int[3][24] ,
         \MR_int[3][23] , \MR_int[3][21] , \MR_int[3][20] , \MR_int[3][19] ,
         \MR_int[3][18] , \MR_int[3][17] , \MR_int[3][16] , \MR_int[3][15] ,
         \MR_int[3][12] , \MR_int[3][11] , \MR_int[3][10] , \MR_int[3][9] ,
         \MR_int[3][8] , \MR_int[3][7] , \MR_int[3][6] , \MR_int[3][4] ,
         \MR_int[3][3] , \MR_int[3][2] , \MR_int[3][1] , \MR_int[4][31] ,
         \MR_int[4][29] , \MR_int[4][28] , \MR_int[4][25] , \MR_int[4][24] ,
         \MR_int[4][22] , \MR_int[4][20] , \MR_int[4][19] , \MR_int[4][18] ,
         \MR_int[4][13] , \MR_int[4][12] , \MR_int[4][11] , \MR_int[4][10] ,
         \MR_int[4][8] , \MR_int[4][6] , \MR_int[4][4] , \MR_int[4][3] ,
         \MR_int[4][2] , \MR_int[5][3] , \MR_int[7][30] , \MR_int[7][29] ,
         \MR_int[7][24] , \MR_int[7][22] , \MR_int[7][20] , \MR_int[7][16] ,
         \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] , \ML_int[1][23] ,
         \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][19] , \ML_int[1][18] ,
         \ML_int[1][17] , \ML_int[1][16] , \ML_int[1][15] , \ML_int[1][14] ,
         \ML_int[1][13] , \ML_int[1][12] , \ML_int[1][11] , \ML_int[1][10] ,
         \ML_int[1][9] , \ML_int[1][8] , \ML_int[1][7] , \ML_int[1][6] ,
         \ML_int[1][5] , \ML_int[1][4] , \ML_int[1][3] , \ML_int[1][2] ,
         \ML_int[1][1] , \ML_int[1][0] , \ML_int[2][31] , \ML_int[2][30] ,
         \ML_int[2][29] , \ML_int[2][28] , \ML_int[2][26] , \ML_int[2][25] ,
         \ML_int[2][24] , \ML_int[2][23] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][17] , \ML_int[2][16] , \ML_int[2][15] ,
         \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] , \ML_int[2][11] ,
         \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] , \ML_int[2][7] ,
         \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] , \ML_int[2][3] ,
         \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] , \ML_int[3][31] ,
         \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] , \ML_int[3][27] ,
         \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] , \ML_int[3][23] ,
         \ML_int[3][21] , \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] ,
         \ML_int[3][16] , \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][15] ,
         \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] , \ML_int[4][11] ,
         \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] , \ML_int[5][31] ,
         \ML_int[5][30] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][18] , \ML_int[5][17] , \ML_int[7][29] , \ML_int[7][28] ,
         \ML_int[7][16] , \ML_int[7][14] , \ML_int[7][10] , \ML_int[7][9] ,
         \ML_int[7][7] , \ML_int[7][6] , \ML_int[7][5] , \ML_int[7][3] ,
         \ML_int[7][2] , \ML_int[7][1] , \ML_int[7][0] , n15, n80, n81, n82,
         n84, n85, n86, n87, n88, n90, n92, n98, n104, net60450, net60477,
         net60578, net60604, net60660, net60751, net60750, net60763, net60869,
         net60893, net61039, net61046, net61053, net61132, net61266, net61331,
         net61353, net61364, net61363, net61624, net61724, net61755, net61774,
         net61783, net61782, net61842, net61851, \ML_int[1][20] ,
         \ML_int[3][22] , \ML_int[2][22] , \ML_int[2][18] , net65464, net65465,
         \temp_int_SH[0] , net61465, n99, n97, n91, n101, n100,
         \MR_int[2][14] , \MR_int[4][30] , \MR_int[1][20] , \MR_int[1][18] ,
         net60718, \ML_int[7][13] , net61436, net60589, net60588,
         \MR_int[4][14] , \MR_int[3][22] , \MR_int[3][14] , \MR_int[2][18] ,
         n121, n122, n124, n125, n131, n132, n135, n136, n138, n139, n141,
         n142, n144, n145, n147, n148, n150, n151, n153, n154, n155, n156,
         n157, n158, n160, n161, n162, n163, n164, n168, n170, n171, n173,
         n174, n175, n178, n180, n181, n182, n183, n184, n186, n189, n192,
         n193, n195, n196, n197, n199, n200, n201, n204, n205, n207, n208,
         n210, n211, n212, n213, n214, n215, n219, n220, n221, n223, n224,
         n225, n226, n227, n228, n229, n230, n232, n233, n234, n235, n236,
         n237, n241, n243, n244, n245, n246, n250, n251, n252, n253, n255,
         n256, n257, n261, n264, n267, n270, n271, n272, n273, n274, n279,
         n282, n283, n284, n285, n286, n295, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n318, n319, n320, n321, n324, n325, n326, n327,
         n328, n329, n331, n332, n333, n334, n335, n336, n337, n338, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n369, n370, n375, n376, n377, n378, n379,
         n380, n381, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n502, n503, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n574, n575, n576,
         n577, n578, n579, n580, n581, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n622, n623, n624, n627, n628, net131991, net134827, net134825,
         net134821, net134819, net134815, net134813, net134811, net134809,
         net134837, net134833, net134831, net134867, net134865, net134861,
         net134859, net134855, net134853, net134851, net134849, net134847,
         net134845, net134843, net134839, net134881, net134879, net134875,
         net134913, net134911, net134905, net134903, net134901, net134899,
         net134897, net134895, net134893, net134891, net134889, net134887,
         net134885, net134883, net134929, net134927, net134925, net134923,
         net134967, net134963, net134959, net134957, net134953, net134951,
         net134949, net134947, net134945, net134943, net134941, net134939,
         net134937, net134935, net134933, net134971, net134969, net134977,
         net134975, net135715, net135717, net135729, net135734, net135859,
         net135858, net135867, net135866, net135876, net135875, net141178,
         net141255, net141408, net141430, net141429, net141428, net141444,
         net141464, net141501, net141507, net141516, net141528, net141534,
         net141544, net141543, net141562, net141563, net141573, n290, n289,
         n288, n287, n109, n108, n107, n106, n96, n89, \MR_int[1][19] ,
         net60313, n292, n291, n110, \temp_int_SH[3] , \temp_int_SH[1] ,
         net60576, net141212, net135865, n95, \MR_int[1][17] ,
         \temp_int_SH[2] , net134965, net134909, n548, n547, n260,
         \MR_int[2][17] , \MR_int[2][13] , net135874, net131988, n83, n340,
         \ML_int[7][4] , net134961, net134873, net134863, \MR_int[3][13] ,
         net134871, net134869, net134841, n128, n127, \MR_int[4][5] ,
         \MR_int[3][5] , n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758;

  MUX2_X1 M1_3_3 ( .A(\MR_int[3][3] ), .B(\MR_int[3][11] ), .S(net134837), .Z(
        \MR_int[4][3] ) );
  MUX2_X1 M1_3_2 ( .A(\MR_int[3][2] ), .B(\MR_int[3][10] ), .S(net134831), .Z(
        \MR_int[4][2] ) );
  MUX2_X1 M1_2_6_0 ( .A(\MR_int[2][6] ), .B(\MR_int[2][10] ), .S(net134929), 
        .Z(\MR_int[3][6] ) );
  MUX2_X1 M1_2_4_0 ( .A(\MR_int[2][4] ), .B(\MR_int[2][8] ), .S(net134927), 
        .Z(\MR_int[3][4] ) );
  MUX2_X1 M1_2_3 ( .A(\MR_int[2][3] ), .B(\MR_int[2][7] ), .S(net134929), .Z(
        \MR_int[3][3] ) );
  MUX2_X1 M1_1_11_0 ( .A(\MR_int[1][11] ), .B(\MR_int[1][13] ), .S(net135859), 
        .Z(\MR_int[2][11] ) );
  MUX2_X1 M1_1_10_0 ( .A(\MR_int[1][10] ), .B(\MR_int[1][12] ), .S(net135858), 
        .Z(\MR_int[2][10] ) );
  MUX2_X1 M1_1_4_0 ( .A(\MR_int[1][4] ), .B(\MR_int[1][6] ), .S(net141464), 
        .Z(\MR_int[2][4] ) );
  MUX2_X1 M1_1_3_0 ( .A(\MR_int[1][3] ), .B(\MR_int[1][5] ), .S(net135859), 
        .Z(\MR_int[2][3] ) );
  MUX2_X1 M1_1_1 ( .A(\MR_int[1][1] ), .B(\ML_int[1][4] ), .S(net141464), .Z(
        \MR_int[2][1] ) );
  MUX2_X1 M1_0_29_0 ( .A(A[29]), .B(A[30]), .S(net141563), .Z(\MR_int[1][29] )
         );
  MUX2_X1 M1_0_28_0 ( .A(A[28]), .B(A[29]), .S(net141408), .Z(\MR_int[1][28] )
         );
  MUX2_X1 M1_0_24_0 ( .A(A[24]), .B(A[25]), .S(net131991), .Z(\MR_int[1][24] )
         );
  MUX2_X1 M1_0_22_0 ( .A(A[22]), .B(A[23]), .S(net141516), .Z(\MR_int[1][22] )
         );
  MUX2_X1 M1_0_9_0 ( .A(A[9]), .B(A[10]), .S(n742), .Z(\MR_int[1][9] ) );
  MUX2_X1 M1_0_8_0 ( .A(A[8]), .B(A[9]), .S(n742), .Z(\MR_int[1][8] ) );
  MUX2_X1 M1_0_6_0 ( .A(A[6]), .B(A[7]), .S(net135729), .Z(\MR_int[1][6] ) );
  MUX2_X1 M1_0_5_0 ( .A(A[5]), .B(A[6]), .S(net141255), .Z(\MR_int[1][5] ) );
  MUX2_X1 M1_0_4_0 ( .A(A[4]), .B(A[5]), .S(n695), .Z(\MR_int[1][4] ) );
  MUX2_X1 M1_0_2_0 ( .A(A[2]), .B(A[3]), .S(net141516), .Z(\MR_int[1][2] ) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(net134811), 
        .Z(\ML_int[5][25] ) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(n755), .S(net134811), .Z(
        \ML_int[5][18] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(net134855), 
        .Z(\ML_int[4][21] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(net134905), 
        .Z(\ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(net134903), 
        .Z(\ML_int[2][30] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(n297), .S(net134903), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(net134901), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n693), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n693), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(net141430), .Z(\ML_int[1][28] )
         );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(net141428), .Z(\ML_int[1][26] )
         );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(net141429), .Z(\ML_int[1][25] )
         );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(net61851), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(net61851), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n705), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n693), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(net141429), .Z(\ML_int[1][14] )
         );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(net135865), .Z(\ML_int[1][13] )
         );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n705), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(net135865), .Z(\ML_int[1][11] )
         );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(net61851), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(net141428), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n710), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(net135866), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(net135865), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(net61851), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(net141430), .Z(\ML_int[1][1] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(net141428), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(net141430), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(net141430), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(net134905), 
        .Z(\ML_int[2][24] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n694), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_13_0 ( .A(A[13]), .B(A[14]), .S(n742), .Z(\MR_int[1][13] ) );
  MUX2_X1 M1_0_1_0 ( .A(A[1]), .B(A[2]), .S(net135729), .Z(\MR_int[1][1] ) );
  MUX2_X1 M1_3_22_0 ( .A(n727), .B(\MR_int[3][30] ), .S(net134837), .Z(
        \MR_int[4][22] ) );
  MUX2_X1 M1_3_11_0 ( .A(\MR_int[3][11] ), .B(\MR_int[3][19] ), .S(net134837), 
        .Z(\MR_int[4][11] ) );
  MUX2_X1 M1_3_14_0 ( .A(n669), .B(n727), .S(net134833), .Z(\MR_int[4][14] )
         );
  MUX2_X1 M1_2_27_0 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(net134923), 
        .Z(\MR_int[3][27] ) );
  MUX2_X1 U3 ( .A(\ML_int[2][26] ), .B(\ML_int[2][30] ), .S(net134923), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 U9 ( .A(\MR_int[2][6] ), .B(\MR_int[2][2] ), .S(net134953), .Z(
        \MR_int[3][2] ) );
  MUX2_X1 U47 ( .A(\ML_int[3][23] ), .B(\ML_int[3][31] ), .S(net134833), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 U78 ( .A(\ML_int[7][16] ), .B(\MR_int[7][16] ), .S(net135876), .Z(
        B[16]) );
  MUX2_X1 U93 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(net134855), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 U127 ( .A(A[22]), .B(A[23]), .S(net141534), .Z(n186) );
  MUX2_X1 U197 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(net134923), .Z(
        n236) );
  MUX2_X1 U204 ( .A(\MR_int[3][10] ), .B(\MR_int[3][18] ), .S(net134837), .Z(
        \MR_int[4][10] ) );
  MUX2_X1 U226 ( .A(\MR_int[2][11] ), .B(\MR_int[2][7] ), .S(net134953), .Z(
        \MR_int[3][7] ) );
  MUX2_X1 U228 ( .A(\MR_int[1][9] ), .B(\MR_int[1][7] ), .S(net134905), .Z(
        \MR_int[2][7] ) );
  MUX2_X1 U235 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(net134903), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 U236 ( .A(\ML_int[2][18] ), .B(\ML_int[2][22] ), .S(net134927), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 U241 ( .A(\ML_int[1][11] ), .B(n728), .S(net134881), .Z(n264) );
  MUX2_X1 U248 ( .A(\ML_int[3][9] ), .B(\ML_int[3][17] ), .S(net134833), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 U254 ( .A(\ML_int[1][24] ), .B(\ML_int[1][26] ), .S(n692), .Z(
        \ML_int[2][26] ) );
  NAND3_X1 U269 ( .A1(\ML_int[5][25] ), .A2(n85), .A3(net134977), .ZN(n336) );
  NAND3_X1 U271 ( .A1(\ML_int[5][24] ), .A2(n85), .A3(net134977), .ZN(n527) );
  MUX2_X1 U288 ( .A(\MR_int[1][20] ), .B(\MR_int[1][18] ), .S(net134903), .Z(
        \MR_int[2][18] ) );
  MUX2_X1 U294 ( .A(\MR_int[3][22] ), .B(\MR_int[3][30] ), .S(net134831), .Z(
        net61774) );
  MUX2_X1 U370 ( .A(\MR_int[3][4] ), .B(\MR_int[3][12] ), .S(net134837), .Z(
        \MR_int[4][4] ) );
  MUX2_X1 U374 ( .A(A[26]), .B(A[25]), .S(n705), .Z(n297) );
  MUX2_X1 U389 ( .A(A[11]), .B(A[10]), .S(n693), .Z(\MR_int[1][10] ) );
  MUX2_X1 U448 ( .A(A[8]), .B(A[7]), .S(net141430), .Z(\MR_int[1][7] ) );
  MUX2_X1 U493 ( .A(A[28]), .B(A[27]), .S(n710), .Z(\MR_int[1][27] ) );
  MUX2_X1 U557 ( .A(A[4]), .B(A[3]), .S(n693), .Z(\MR_int[1][3] ) );
  MUX2_X1 U558 ( .A(A[30]), .B(A[31]), .S(net141212), .Z(\MR_int[1][30] ) );
  MUX2_X1 U565 ( .A(A[13]), .B(A[12]), .S(net141429), .Z(\MR_int[1][12] ) );
  MUX2_X1 U601 ( .A(\MR_int[1][12] ), .B(\MR_int[1][14] ), .S(net135858), .Z(
        n410) );
  MUX2_X1 U621 ( .A(A[27]), .B(A[26]), .S(net141429), .Z(n424) );
  MUX2_X1 U734 ( .A(A[16]), .B(A[15]), .S(n694), .Z(\MR_int[1][15] ) );
  MUX2_X1 U768 ( .A(A[15]), .B(A[14]), .S(n729), .Z(\MR_int[1][14] ) );
  MUX2_X1 U777 ( .A(\MR_int[3][16] ), .B(\MR_int[3][8] ), .S(net134855), .Z(
        \MR_int[4][8] ) );
  MUX2_X1 U913 ( .A(A[23]), .B(A[24]), .S(n742), .Z(n601) );
  MUX2_X1 U299 ( .A(n424), .B(\ML_int[1][25] ), .S(net134901), .Z(n250) );
  MUX2_X1 U732 ( .A(\ML_int[7][29] ), .B(\MR_int[7][29] ), .S(net135876), .Z(
        B[29]) );
  AND2_X2 U273 ( .A1(\SHMAG[5] ), .A2(net134977), .ZN(n85) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(net134953), .Z(
        \ML_int[3][4] ) );
  NAND3_X1 U365 ( .A1(SH[16]), .A2(SH[15]), .A3(SH[14]), .ZN(net60751) );
  NAND3_X1 U364 ( .A1(SH[18]), .A2(SH[17]), .A3(SH[19]), .ZN(net61363) );
  NAND3_X1 U281 ( .A1(SH[22]), .A2(SH[21]), .A3(SH[20]), .ZN(net61364) );
  MUX2_X1 M1_0_20_0 ( .A(A[20]), .B(A[21]), .S(net141408), .Z(\MR_int[1][20] )
         );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(net61851), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n710), .Z(\ML_int[1][21] ) );
  NAND3_X1 U367 ( .A1(SH[8]), .A2(SH[7]), .A3(SH[9]), .ZN(net65464) );
  NAND3_X1 U368 ( .A1(SH[30]), .A2(SH[29]), .A3(SH[6]), .ZN(net65465) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(net61851), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(net141429), .Z(\ML_int[1][17] )
         );
  MUX2_X1 M1_0_16_0 ( .A(A[16]), .B(A[17]), .S(net141563), .Z(\MR_int[1][16] )
         );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(net141544), .Z(\ML_int[1][18] )
         );
  MUX2_X1 M1_0_25_0 ( .A(A[25]), .B(A[26]), .S(net141212), .Z(\MR_int[1][25] )
         );
  MUX2_X1 M1_0_17_0 ( .A(A[17]), .B(A[18]), .S(net141178), .Z(\MR_int[1][17] )
         );
  MUX2_X1 M1_2_5_0 ( .A(\MR_int[2][5] ), .B(\MR_int[2][9] ), .S(net134925), 
        .Z(\MR_int[3][5] ) );
  NAND4_X1 U4 ( .A1(n109), .A2(n110), .A3(n107), .A4(n108), .ZN(n656) );
  BUF_X1 U5 ( .A(\temp_int_SH[0] ), .Z(net135865) );
  AND3_X1 U6 ( .A1(n657), .A2(n658), .A3(n659), .ZN(n109) );
  NOR2_X1 U7 ( .A1(SH[27]), .A2(SH[26]), .ZN(n657) );
  AND2_X1 U8 ( .A1(n721), .A2(n719), .ZN(n658) );
  AND2_X1 U10 ( .A1(n720), .A2(n718), .ZN(n659) );
  BUF_X1 U11 ( .A(net134961), .Z(net134939) );
  NAND2_X1 U12 ( .A1(\MR_int[3][26] ), .A2(net134833), .ZN(n660) );
  INV_X1 U13 ( .A(net141501), .ZN(net141429) );
  INV_X2 U14 ( .A(net134967), .ZN(net134925) );
  NAND2_X1 U15 ( .A1(\MR_int[3][17] ), .A2(n664), .ZN(n661) );
  NAND2_X1 U16 ( .A1(n661), .A2(n662), .ZN(\MR_int[7][16] ) );
  OR2_X1 U17 ( .A1(n663), .A2(n243), .ZN(n662) );
  INV_X1 U18 ( .A(n205), .ZN(n663) );
  AND2_X1 U19 ( .A1(net134839), .A2(n205), .ZN(n664) );
  CLKBUF_X1 U20 ( .A(n579), .Z(n665) );
  BUF_X2 U21 ( .A(net134911), .Z(net134897) );
  NAND2_X1 U22 ( .A1(n723), .A2(n666), .ZN(B[11]) );
  AND2_X1 U23 ( .A1(n724), .A2(n532), .ZN(n666) );
  INV_X2 U24 ( .A(net141501), .ZN(net141430) );
  NAND2_X1 U25 ( .A1(\MR_int[4][14] ), .A2(n170), .ZN(n667) );
  NAND2_X1 U26 ( .A1(n667), .A2(n668), .ZN(B[13]) );
  AND2_X1 U27 ( .A1(net60718), .A2(n168), .ZN(n668) );
  NAND2_X1 U28 ( .A1(net60588), .A2(net60589), .ZN(n669) );
  MUX2_X1 U29 ( .A(A[30]), .B(A[29]), .S(net135867), .Z(\ML_int[1][30] ) );
  CLKBUF_X1 U30 ( .A(n689), .Z(n670) );
  BUF_X1 U31 ( .A(\temp_int_SH[2] ), .Z(net134967) );
  INV_X1 U32 ( .A(net134965), .ZN(net134929) );
  BUF_X1 U33 ( .A(net134911), .Z(net134883) );
  INV_X1 U34 ( .A(\temp_int_SH[2] ), .ZN(net134927) );
  INV_X1 U35 ( .A(net134827), .ZN(net134811) );
  BUF_X1 U36 ( .A(net134911), .Z(net134903) );
  NAND2_X1 U37 ( .A1(net134927), .A2(net134865), .ZN(n671) );
  NAND2_X1 U38 ( .A1(n85), .A2(net134977), .ZN(n672) );
  NAND2_X1 U39 ( .A1(\MR_int[3][1] ), .A2(net134855), .ZN(n673) );
  BUF_X1 U40 ( .A(SH[31]), .Z(net135875) );
  BUF_X1 U41 ( .A(net131988), .Z(net134975) );
  MUX2_X1 U42 ( .A(\MR_int[3][12] ), .B(\MR_int[3][20] ), .S(net134837), .Z(
        \MR_int[4][12] ) );
  CLKBUF_X1 U43 ( .A(SH[31]), .Z(net135874) );
  MUX2_X1 U44 ( .A(\MR_int[1][13] ), .B(\MR_int[1][15] ), .S(net134881), .Z(
        \MR_int[2][13] ) );
  BUF_X1 U45 ( .A(\temp_int_SH[1] ), .Z(net134909) );
  MUX2_X1 U46 ( .A(A[19]), .B(A[18]), .S(net141544), .Z(\MR_int[1][18] ) );
  BUF_X1 U48 ( .A(SH[31]), .Z(net135876) );
  AND2_X1 U49 ( .A1(n303), .A2(n304), .ZN(n674) );
  NOR2_X1 U50 ( .A1(n675), .A2(n676), .ZN(n679) );
  AND2_X1 U51 ( .A1(n606), .A2(n607), .ZN(n675) );
  NAND2_X1 U52 ( .A1(net134971), .A2(n716), .ZN(n676) );
  OAI21_X1 U53 ( .B1(n678), .B2(n679), .A(net135875), .ZN(n677) );
  AND2_X1 U54 ( .A1(\MR_int[4][5] ), .A2(n205), .ZN(n678) );
  OAI21_X1 U55 ( .B1(net134925), .B2(n680), .A(n503), .ZN(\ML_int[3][19] ) );
  INV_X1 U56 ( .A(\ML_int[2][15] ), .ZN(n680) );
  OAI221_X1 U57 ( .B1(n681), .B2(n476), .C1(n224), .C2(n737), .A(n502), .ZN(
        B[0]) );
  INV_X1 U58 ( .A(n295), .ZN(n681) );
  AOI22_X1 U59 ( .A1(n731), .A2(\ML_int[1][21] ), .B1(n682), .B2(net134923), 
        .ZN(n510) );
  INV_X1 U60 ( .A(n459), .ZN(n682) );
  NAND3_X1 U61 ( .A1(n422), .A2(n225), .A3(n423), .ZN(n163) );
  NAND2_X1 U62 ( .A1(n344), .A2(n343), .ZN(\ML_int[2][15] ) );
  OAI21_X1 U63 ( .B1(n683), .B2(n670), .A(net134833), .ZN(n468) );
  INV_X1 U64 ( .A(n565), .ZN(n683) );
  OAI21_X1 U65 ( .B1(n674), .B2(n672), .A(n572), .ZN(B[19]) );
  OAI21_X1 U66 ( .B1(net134827), .B2(n673), .A(n744), .ZN(n295) );
  MUX2_X1 U67 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(\temp_int_SH[2] ), 
        .Z(\ML_int[3][26] ) );
  AOI21_X1 U68 ( .B1(n193), .B2(n192), .A(net134825), .ZN(n684) );
  INV_X1 U69 ( .A(n684), .ZN(n533) );
  AOI21_X1 U70 ( .B1(n702), .B2(n701), .A(n685), .ZN(n686) );
  INV_X1 U71 ( .A(n493), .ZN(n685) );
  INV_X1 U72 ( .A(n686), .ZN(n402) );
  NAND2_X1 U73 ( .A1(n299), .A2(n298), .ZN(\ML_int[5][26] ) );
  NAND3_X1 U74 ( .A1(n232), .A2(n233), .A3(n594), .ZN(B[9]) );
  NAND2_X1 U75 ( .A1(net134879), .A2(\MR_int[1][14] ), .ZN(n343) );
  INV_X2 U76 ( .A(net134911), .ZN(net134879) );
  OAI22_X1 U77 ( .A1(n687), .A2(n671), .B1(net61039), .B2(net134837), .ZN(n688) );
  INV_X1 U79 ( .A(n348), .ZN(n687) );
  INV_X1 U80 ( .A(n688), .ZN(n489) );
  NAND3_X1 U81 ( .A1(n363), .A2(n409), .A3(n364), .ZN(\ML_int[4][9] ) );
  AOI21_X1 U82 ( .B1(n547), .B2(n548), .A(net134923), .ZN(n689) );
  INV_X1 U83 ( .A(n689), .ZN(n564) );
  AOI21_X1 U84 ( .B1(n468), .B2(n467), .A(net134825), .ZN(n690) );
  INV_X1 U85 ( .A(n690), .ZN(n411) );
  AOI21_X1 U86 ( .B1(n589), .B2(n588), .A(n476), .ZN(n691) );
  INV_X1 U87 ( .A(n691), .ZN(n610) );
  INV_X1 U88 ( .A(net134905), .ZN(n692) );
  BUF_X2 U89 ( .A(net134909), .Z(net134905) );
  BUF_X1 U90 ( .A(net135734), .Z(n693) );
  BUF_X1 U91 ( .A(n729), .Z(n694) );
  BUF_X1 U92 ( .A(\temp_int_SH[0] ), .Z(net141544) );
  BUF_X1 U94 ( .A(net134913), .Z(net134901) );
  BUF_X1 U95 ( .A(net134967), .Z(net134959) );
  MUX2_X1 U96 ( .A(\MR_int[1][20] ), .B(\MR_int[1][18] ), .S(net134897), .Z(
        net61353) );
  INV_X1 U97 ( .A(net141544), .ZN(n695) );
  AND2_X1 U98 ( .A1(n583), .A2(n213), .ZN(n696) );
  NAND2_X1 U99 ( .A1(\ML_int[4][22] ), .A2(net134815), .ZN(n697) );
  NAND2_X1 U100 ( .A1(n752), .A2(net134811), .ZN(n698) );
  NAND2_X1 U101 ( .A1(n697), .A2(n698), .ZN(\ML_int[5][22] ) );
  CLKBUF_X1 U102 ( .A(net134913), .Z(net134887) );
  CLKBUF_X1 U103 ( .A(net134911), .Z(net134885) );
  NAND2_X1 U104 ( .A1(\ML_int[1][5] ), .A2(net135859), .ZN(n699) );
  NAND2_X1 U105 ( .A1(\ML_int[1][3] ), .A2(net134903), .ZN(n700) );
  NAND2_X1 U106 ( .A1(n699), .A2(n700), .ZN(\ML_int[2][5] ) );
  AND2_X2 U107 ( .A1(n96), .A2(n89), .ZN(net141501) );
  NAND2_X1 U108 ( .A1(\ML_int[4][11] ), .A2(net134813), .ZN(n701) );
  NAND2_X1 U109 ( .A1(\ML_int[4][27] ), .A2(net134815), .ZN(n702) );
  BUF_X1 U110 ( .A(\temp_int_SH[0] ), .Z(net141543) );
  NAND2_X1 U111 ( .A1(\MR_int[4][24] ), .A2(net134811), .ZN(n703) );
  OR2_X1 U112 ( .A1(n703), .A2(n704), .ZN(n515) );
  OR2_X1 U113 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(n704) );
  BUF_X1 U114 ( .A(net135734), .Z(n705) );
  NAND2_X1 U115 ( .A1(\MR_int[1][25] ), .A2(net134879), .ZN(n706) );
  NAND2_X1 U116 ( .A1(n601), .A2(net134903), .ZN(n707) );
  NAND2_X1 U117 ( .A1(n706), .A2(n707), .ZN(\MR_int[2][23] ) );
  AND2_X1 U118 ( .A1(n708), .A2(n709), .ZN(n446) );
  NAND2_X1 U119 ( .A1(\MR_int[4][13] ), .A2(n204), .ZN(n708) );
  OR2_X1 U120 ( .A1(n359), .A2(n456), .ZN(n709) );
  BUF_X1 U121 ( .A(net135734), .Z(n710) );
  NAND2_X1 U122 ( .A1(\ML_int[1][30] ), .A2(n711), .ZN(n712) );
  NAND2_X1 U123 ( .A1(\MR_int[1][27] ), .A2(net134901), .ZN(n713) );
  NAND2_X1 U124 ( .A1(n712), .A2(n713), .ZN(\MR_int[2][27] ) );
  INV_X1 U125 ( .A(net134901), .ZN(n711) );
  NAND2_X1 U126 ( .A1(\ML_int[4][30] ), .A2(net134815), .ZN(n714) );
  NAND2_X1 U128 ( .A1(\ML_int[4][14] ), .A2(net134811), .ZN(n715) );
  NAND2_X1 U129 ( .A1(n714), .A2(n715), .ZN(\ML_int[5][30] ) );
  INV_X1 U130 ( .A(\SHMAG[5] ), .ZN(n716) );
  AND2_X1 U131 ( .A1(net134813), .A2(n716), .ZN(n205) );
  NAND2_X1 U132 ( .A1(n716), .A2(n274), .ZN(n271) );
  BUF_X2 U133 ( .A(n173), .Z(net134971) );
  NAND2_X1 U134 ( .A1(n127), .A2(n128), .ZN(\MR_int[4][5] ) );
  NAND2_X1 U135 ( .A1(\MR_int[3][5] ), .A2(net134841), .ZN(n128) );
  BUF_X1 U136 ( .A(net134869), .Z(net134841) );
  NAND2_X1 U137 ( .A1(\ML_int[3][0] ), .A2(net134841), .ZN(n491) );
  NAND2_X1 U138 ( .A1(\MR_int[3][21] ), .A2(net134841), .ZN(n606) );
  NAND2_X1 U139 ( .A1(\ML_int[3][18] ), .A2(net134841), .ZN(n145) );
  BUF_X1 U140 ( .A(net134871), .Z(net134869) );
  BUF_X1 U141 ( .A(net134869), .Z(net134839) );
  BUF_X1 U142 ( .A(net134869), .Z(net134843) );
  AND2_X1 U143 ( .A1(net134971), .A2(net134869), .ZN(n220) );
  CLKBUF_X1 U144 ( .A(\temp_int_SH[3] ), .Z(net134871) );
  CLKBUF_X1 U145 ( .A(net134871), .Z(net134867) );
  INV_X1 U146 ( .A(net134871), .ZN(net134837) );
  NAND2_X1 U147 ( .A1(\MR_int[3][13] ), .A2(net134833), .ZN(n127) );
  INV_X2 U148 ( .A(net134859), .ZN(net134833) );
  BUF_X2 U149 ( .A(net134863), .Z(net134859) );
  BUF_X1 U150 ( .A(net134873), .Z(net134863) );
  CLKBUF_X1 U151 ( .A(net134863), .Z(net134861) );
  BUF_X1 U152 ( .A(\temp_int_SH[3] ), .Z(net134873) );
  BUF_X1 U153 ( .A(net134873), .Z(net134865) );
  MUX2_X1 U154 ( .A(\MR_int[2][17] ), .B(\MR_int[2][13] ), .S(net134939), .Z(
        \MR_int[3][13] ) );
  BUF_X1 U155 ( .A(net134965), .Z(net134961) );
  BUF_X1 U156 ( .A(net134961), .Z(net134941) );
  BUF_X1 U157 ( .A(net134961), .Z(net134943) );
  BUF_X1 U158 ( .A(\temp_int_SH[2] ), .Z(net134965) );
  NAND2_X1 U159 ( .A1(n677), .A2(n340), .ZN(B[4]) );
  NAND2_X1 U160 ( .A1(\ML_int[7][4] ), .A2(net134977), .ZN(n340) );
  BUF_X4 U161 ( .A(net131988), .Z(net134977) );
  INV_X1 U162 ( .A(net135874), .ZN(net131988) );
  NAND2_X1 U163 ( .A1(n106), .A2(net131988), .ZN(net61465) );
  NAND2_X1 U164 ( .A1(n656), .A2(net131988), .ZN(n89) );
  NOR2_X1 U165 ( .A1(n325), .A2(n83), .ZN(\ML_int[7][4] ) );
  NAND2_X1 U166 ( .A1(net141573), .A2(net134833), .ZN(n83) );
  BUF_X1 U167 ( .A(net134965), .Z(net134963) );
  NAND2_X1 U168 ( .A1(n547), .A2(n548), .ZN(\MR_int[2][17] ) );
  MUX2_X1 U169 ( .A(\MR_int[2][13] ), .B(\MR_int[2][17] ), .S(net134929), .Z(
        net141562) );
  NAND2_X1 U170 ( .A1(\MR_int[1][19] ), .A2(net134875), .ZN(n548) );
  INV_X1 U171 ( .A(net134905), .ZN(net134875) );
  INV_X1 U172 ( .A(net134909), .ZN(net135717) );
  NAND2_X1 U173 ( .A1(\MR_int[1][17] ), .A2(net134897), .ZN(n547) );
  BUF_X2 U174 ( .A(\temp_int_SH[1] ), .Z(net134911) );
  NAND2_X1 U175 ( .A1(\MR_int[2][13] ), .A2(net134927), .ZN(n557) );
  NAND2_X1 U176 ( .A1(net61465), .A2(n260), .ZN(\temp_int_SH[2] ) );
  INV_X1 U177 ( .A(\temp_int_SH[2] ), .ZN(net134923) );
  NAND2_X1 U178 ( .A1(SH[2]), .A2(net141507), .ZN(n260) );
  NAND2_X1 U179 ( .A1(\MR_int[1][19] ), .A2(net134891), .ZN(n595) );
  CLKBUF_X1 U180 ( .A(\temp_int_SH[1] ), .Z(net134913) );
  NAND2_X1 U181 ( .A1(\MR_int[1][17] ), .A2(net134879), .ZN(n581) );
  INV_X1 U182 ( .A(net135867), .ZN(net141212) );
  INV_X1 U183 ( .A(net135867), .ZN(net131991) );
  NAND2_X1 U184 ( .A1(n89), .A2(n95), .ZN(\temp_int_SH[1] ) );
  NAND2_X1 U185 ( .A1(SH[1]), .A2(net60576), .ZN(n95) );
  NAND2_X1 U186 ( .A1(net60578), .A2(net135875), .ZN(net60576) );
  NAND2_X1 U187 ( .A1(n89), .A2(n96), .ZN(\temp_int_SH[0] ) );
  CLKBUF_X1 U188 ( .A(net61465), .Z(net135715) );
  NAND2_X1 U189 ( .A1(net60578), .A2(net135875), .ZN(net141507) );
  NAND2_X1 U190 ( .A1(net61465), .A2(n717), .ZN(\temp_int_SH[3] ) );
  NAND2_X1 U191 ( .A1(SH[3]), .A2(net141507), .ZN(n717) );
  AND3_X1 U192 ( .A1(net60313), .A2(n292), .A3(n291), .ZN(n110) );
  NAND4_X1 U193 ( .A1(n109), .A2(n110), .A3(n107), .A4(n108), .ZN(n106) );
  NOR2_X1 U194 ( .A1(SH[6]), .A2(SH[9]), .ZN(n291) );
  NOR2_X1 U195 ( .A1(SH[8]), .A2(SH[7]), .ZN(n292) );
  NOR3_X1 U196 ( .A1(SH[28]), .A2(SH[29]), .A3(SH[30]), .ZN(net60313) );
  AND3_X1 U198 ( .A1(SH[28]), .A2(SH[26]), .A3(SH[27]), .ZN(net60450) );
  MUX2_X1 U199 ( .A(A[20]), .B(A[19]), .S(net141430), .Z(\MR_int[1][19] ) );
  NAND2_X1 U200 ( .A1(n91), .A2(SH[0]), .ZN(n96) );
  NAND2_X1 U201 ( .A1(n91), .A2(SH[0]), .ZN(net141444) );
  AND2_X1 U202 ( .A1(n287), .A2(n289), .ZN(n108) );
  NOR3_X1 U203 ( .A1(SH[20]), .A2(SH[21]), .A3(SH[19]), .ZN(n289) );
  NOR3_X1 U205 ( .A1(SH[17]), .A2(SH[18]), .A3(SH[16]), .ZN(n287) );
  AND2_X1 U206 ( .A1(n290), .A2(n288), .ZN(n107) );
  NOR3_X1 U207 ( .A1(SH[11]), .A2(SH[12]), .A3(SH[10]), .ZN(n288) );
  NOR3_X1 U208 ( .A1(SH[14]), .A2(SH[15]), .A3(SH[13]), .ZN(n290) );
  INV_X1 U209 ( .A(SH[22]), .ZN(n718) );
  INV_X1 U210 ( .A(SH[24]), .ZN(n720) );
  INV_X1 U211 ( .A(SH[23]), .ZN(n719) );
  INV_X1 U212 ( .A(SH[25]), .ZN(n721) );
  NAND4_X1 U213 ( .A1(SH[11]), .A2(SH[12]), .A3(SH[13]), .A4(SH[10]), .ZN(
        net60750) );
  AND3_X1 U214 ( .A1(SH[24]), .A2(SH[25]), .A3(SH[23]), .ZN(n104) );
  NAND2_X1 U215 ( .A1(\ML_int[2][13] ), .A2(n722), .ZN(n356) );
  AND2_X1 U216 ( .A1(net134929), .A2(net134837), .ZN(n722) );
  MUX2_X1 U217 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(net134953), .Z(
        net141573) );
  NAND2_X1 U218 ( .A1(\MR_int[4][12] ), .A2(n241), .ZN(n723) );
  OR2_X1 U219 ( .A1(n208), .A2(n592), .ZN(n724) );
  BUF_X1 U220 ( .A(\temp_int_SH[0] ), .Z(net135866) );
  MUX2_X1 U221 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(net134925), .Z(
        n725) );
  MUX2_X1 U222 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(net134923), .Z(
        n726) );
  NAND2_X1 U223 ( .A1(n279), .A2(net60477), .ZN(n727) );
  INV_X1 U224 ( .A(net135866), .ZN(net141563) );
  MUX2_X1 U225 ( .A(A[13]), .B(A[12]), .S(net141544), .Z(n728) );
  MUX2_X1 U227 ( .A(A[27]), .B(A[26]), .S(net141429), .Z(\MR_int[1][26] ) );
  INV_X1 U229 ( .A(net141428), .ZN(net141534) );
  INV_X1 U230 ( .A(net134905), .ZN(net141528) );
  INV_X1 U231 ( .A(net141428), .ZN(net141516) );
  NAND2_X1 U232 ( .A1(net61465), .A2(net141444), .ZN(n729) );
  NAND2_X1 U233 ( .A1(net61465), .A2(net141444), .ZN(net61851) );
  INV_X1 U234 ( .A(net134897), .ZN(net141464) );
  BUF_X2 U237 ( .A(net135717), .Z(net135858) );
  INV_X1 U238 ( .A(net141501), .ZN(net141428) );
  INV_X1 U239 ( .A(net141543), .ZN(net141408) );
  NAND2_X1 U240 ( .A1(n484), .A2(n485), .ZN(n730) );
  AND2_X1 U242 ( .A1(net135858), .A2(net134927), .ZN(n731) );
  MUX2_X1 U243 ( .A(A[12]), .B(A[11]), .S(net141430), .Z(\MR_int[1][11] ) );
  MUX2_X1 U244 ( .A(A[28]), .B(A[29]), .S(net141534), .Z(n732) );
  NAND2_X1 U245 ( .A1(\ML_int[4][29] ), .A2(n733), .ZN(n735) );
  NOR2_X1 U246 ( .A1(n758), .A2(net134813), .ZN(n733) );
  MUX2_X2 U247 ( .A(\MR_int[2][30] ), .B(\MR_int[2][26] ), .S(net134967), .Z(
        \MR_int[3][26] ) );
  NAND2_X1 U249 ( .A1(\ML_int[4][13] ), .A2(n736), .ZN(n734) );
  NAND2_X1 U250 ( .A1(n735), .A2(n734), .ZN(\ML_int[7][29] ) );
  AND2_X1 U251 ( .A1(net134809), .A2(n85), .ZN(n736) );
  INV_X1 U252 ( .A(net141543), .ZN(net135729) );
  INV_X1 U253 ( .A(net135866), .ZN(net141255) );
  OR2_X1 U255 ( .A1(net134811), .A2(n476), .ZN(n737) );
  BUF_X2 U256 ( .A(net134957), .Z(net134953) );
  BUF_X1 U257 ( .A(net134957), .Z(net134951) );
  CLKBUF_X1 U258 ( .A(net134911), .Z(net134889) );
  INV_X1 U259 ( .A(net141543), .ZN(net141178) );
  INV_X1 U260 ( .A(n88), .ZN(n757) );
  INV_X1 U261 ( .A(n87), .ZN(n756) );
  NAND2_X1 U262 ( .A1(n753), .A2(net134809), .ZN(n125) );
  INV_X1 U263 ( .A(n82), .ZN(n753) );
  OR2_X1 U264 ( .A1(net134811), .A2(n603), .ZN(n183) );
  INV_X1 U265 ( .A(n84), .ZN(n754) );
  INV_X1 U266 ( .A(net134825), .ZN(net134809) );
  AND2_X1 U267 ( .A1(n477), .A2(n256), .ZN(n178) );
  INV_X1 U268 ( .A(net134905), .ZN(net134881) );
  NOR2_X1 U270 ( .A1(n325), .A2(n84), .ZN(\ML_int[7][3] ) );
  NOR2_X1 U272 ( .A1(n325), .A2(n81), .ZN(\ML_int[7][6] ) );
  BUF_X1 U274 ( .A(net134865), .Z(net134855) );
  BUF_X1 U275 ( .A(net134867), .Z(net134847) );
  NOR2_X1 U276 ( .A1(net134925), .A2(n751), .ZN(\MR_int[3][30] ) );
  NAND2_X1 U277 ( .A1(\ML_int[3][3] ), .A2(net134833), .ZN(n84) );
  NAND2_X1 U278 ( .A1(\ML_int[3][2] ), .A2(net134833), .ZN(n86) );
  CLKBUF_X1 U279 ( .A(net134865), .Z(net134853) );
  BUF_X1 U280 ( .A(net134963), .Z(net134935) );
  BUF_X1 U282 ( .A(net134963), .Z(net134933) );
  BUF_X1 U283 ( .A(net134867), .Z(net134845) );
  BUF_X1 U284 ( .A(net134959), .Z(net134945) );
  BUF_X1 U285 ( .A(net134867), .Z(net134849) );
  NAND2_X1 U286 ( .A1(\ML_int[3][14] ), .A2(net134831), .ZN(n550) );
  NAND2_X1 U287 ( .A1(\ML_int[3][6] ), .A2(net134851), .ZN(n551) );
  NAND2_X1 U289 ( .A1(n174), .A2(net134833), .ZN(n423) );
  NAND2_X1 U290 ( .A1(n445), .A2(n444), .ZN(n174) );
  BUF_X1 U291 ( .A(net134865), .Z(net134851) );
  NAND2_X1 U292 ( .A1(n416), .A2(n415), .ZN(\ML_int[4][12] ) );
  BUF_X1 U293 ( .A(net134963), .Z(net134937) );
  BUF_X1 U295 ( .A(net134959), .Z(net134949) );
  NAND2_X1 U296 ( .A1(n437), .A2(n438), .ZN(\ML_int[4][11] ) );
  NAND2_X1 U297 ( .A1(\ML_int[3][3] ), .A2(net134847), .ZN(n438) );
  NAND2_X1 U298 ( .A1(\ML_int[3][11] ), .A2(net134837), .ZN(n437) );
  NAND2_X1 U300 ( .A1(n400), .A2(n399), .ZN(\ML_int[4][20] ) );
  NAND2_X1 U301 ( .A1(n253), .A2(net134831), .ZN(n399) );
  NAND2_X1 U302 ( .A1(net61132), .A2(n475), .ZN(\ML_int[4][15] ) );
  NAND2_X1 U303 ( .A1(\ML_int[3][7] ), .A2(net134847), .ZN(n475) );
  NAND2_X1 U304 ( .A1(\ML_int[3][15] ), .A2(net134831), .ZN(net61132) );
  NAND2_X1 U305 ( .A1(\ML_int[4][8] ), .A2(n622), .ZN(n267) );
  NAND2_X1 U306 ( .A1(n490), .A2(n491), .ZN(\ML_int[4][8] ) );
  NAND2_X1 U307 ( .A1(\ML_int[3][8] ), .A2(net134831), .ZN(n490) );
  BUF_X1 U308 ( .A(net134959), .Z(net134947) );
  NAND2_X1 U309 ( .A1(\ML_int[3][16] ), .A2(net134853), .ZN(n432) );
  NAND2_X1 U310 ( .A1(\ML_int[4][19] ), .A2(net134819), .ZN(n303) );
  NAND2_X1 U311 ( .A1(\ML_int[3][11] ), .A2(net134845), .ZN(n426) );
  NAND2_X1 U312 ( .A1(n138), .A2(n139), .ZN(\ML_int[4][10] ) );
  NAND2_X1 U313 ( .A1(\ML_int[3][2] ), .A2(net134847), .ZN(n139) );
  NAND2_X1 U314 ( .A1(\ML_int[5][17] ), .A2(n379), .ZN(n450) );
  NAND2_X1 U315 ( .A1(n360), .A2(n361), .ZN(\ML_int[5][17] ) );
  NAND2_X1 U316 ( .A1(n756), .A2(net134809), .ZN(n361) );
  AND2_X1 U317 ( .A1(net134861), .A2(net134971), .ZN(n184) );
  NAND2_X1 U318 ( .A1(\ML_int[5][20] ), .A2(n227), .ZN(n443) );
  NAND2_X1 U319 ( .A1(n366), .A2(n367), .ZN(\ML_int[5][20] ) );
  NAND2_X1 U320 ( .A1(n309), .A2(net134809), .ZN(n367) );
  NAND2_X1 U321 ( .A1(\ML_int[4][20] ), .A2(net134819), .ZN(n366) );
  NAND2_X1 U322 ( .A1(n513), .A2(n512), .ZN(\ML_int[4][23] ) );
  NAND2_X1 U323 ( .A1(\ML_int[3][23] ), .A2(net134831), .ZN(n513) );
  NAND2_X1 U324 ( .A1(\ML_int[3][15] ), .A2(net134845), .ZN(n512) );
  NAND2_X1 U325 ( .A1(\ML_int[3][22] ), .A2(net134847), .ZN(net61053) );
  AND2_X1 U326 ( .A1(\ML_int[3][16] ), .A2(n158), .ZN(n161) );
  AND2_X1 U327 ( .A1(\ML_int[3][8] ), .A2(n199), .ZN(n160) );
  AND2_X1 U328 ( .A1(net134861), .A2(n252), .ZN(n199) );
  AND2_X1 U329 ( .A1(\ML_int[4][9] ), .A2(n622), .ZN(\ML_int[7][9] ) );
  NAND2_X1 U330 ( .A1(\ML_int[3][8] ), .A2(n246), .ZN(n244) );
  OR2_X1 U331 ( .A1(n197), .A2(net134971), .ZN(n388) );
  OR2_X1 U332 ( .A1(n750), .A2(net134971), .ZN(n324) );
  INV_X1 U333 ( .A(\MR_int[4][28] ), .ZN(n750) );
  OR2_X1 U334 ( .A1(net134825), .A2(n491), .ZN(n245) );
  NAND2_X1 U335 ( .A1(\ML_int[5][23] ), .A2(n379), .ZN(n514) );
  NAND2_X1 U336 ( .A1(n471), .A2(n472), .ZN(\ML_int[5][23] ) );
  OR2_X1 U337 ( .A1(n80), .A2(net134827), .ZN(n472) );
  NAND2_X1 U338 ( .A1(\ML_int[4][23] ), .A2(net134819), .ZN(n471) );
  OR2_X1 U339 ( .A1(n466), .A2(net134859), .ZN(n364) );
  NAND2_X1 U340 ( .A1(n470), .A2(n469), .ZN(\ML_int[5][24] ) );
  NAND2_X1 U341 ( .A1(\ML_int[4][24] ), .A2(net134969), .ZN(n470) );
  AND2_X1 U342 ( .A1(n244), .A2(n245), .ZN(n469) );
  NAND2_X1 U343 ( .A1(n431), .A2(n432), .ZN(\ML_int[4][24] ) );
  INV_X1 U344 ( .A(n86), .ZN(n755) );
  NAND2_X1 U345 ( .A1(n369), .A2(n370), .ZN(\ML_int[4][18] ) );
  NAND2_X1 U346 ( .A1(n430), .A2(n429), .ZN(\ML_int[4][27] ) );
  NAND2_X1 U347 ( .A1(n328), .A2(n329), .ZN(\ML_int[7][16] ) );
  OR2_X1 U348 ( .A1(n758), .A2(n362), .ZN(n329) );
  NOR2_X1 U349 ( .A1(n160), .A2(n161), .ZN(n328) );
  NAND2_X1 U350 ( .A1(n757), .A2(net134811), .ZN(n362) );
  AND2_X1 U351 ( .A1(\ML_int[4][10] ), .A2(n622), .ZN(\ML_int[7][10] ) );
  NAND2_X1 U352 ( .A1(\ML_int[5][22] ), .A2(n493), .ZN(n495) );
  INV_X1 U353 ( .A(n81), .ZN(n752) );
  INV_X1 U354 ( .A(n225), .ZN(n746) );
  NAND2_X1 U355 ( .A1(n85), .A2(net134969), .ZN(n325) );
  AND2_X1 U356 ( .A1(n85), .A2(net134971), .ZN(n622) );
  NAND2_X1 U357 ( .A1(\ML_int[7][9] ), .A2(net134975), .ZN(n594) );
  NAND2_X1 U358 ( .A1(\ML_int[4][11] ), .A2(n211), .ZN(n532) );
  NAND2_X1 U359 ( .A1(n455), .A2(n454), .ZN(B[15]) );
  NAND2_X1 U360 ( .A1(n384), .A2(n622), .ZN(n455) );
  NAND2_X1 U361 ( .A1(n446), .A2(n447), .ZN(B[12]) );
  NAND2_X1 U362 ( .A1(n235), .A2(n622), .ZN(n447) );
  BUF_X1 U363 ( .A(n173), .Z(net134969) );
  AND2_X1 U366 ( .A1(\ML_int[5][31] ), .A2(n378), .ZN(B[31]) );
  AND2_X1 U369 ( .A1(n85), .A2(net134977), .ZN(n378) );
  AND2_X1 U371 ( .A1(net134813), .A2(n405), .ZN(n383) );
  NAND2_X1 U372 ( .A1(n402), .A2(n401), .ZN(B[27]) );
  OR2_X1 U373 ( .A1(n324), .A2(n359), .ZN(n401) );
  NAND2_X1 U375 ( .A1(\ML_int[7][13] ), .A2(net134975), .ZN(net60718) );
  NAND2_X1 U376 ( .A1(\ML_int[2][6] ), .A2(net134927), .ZN(n586) );
  NAND2_X1 U377 ( .A1(\ML_int[2][2] ), .A2(net134941), .ZN(n587) );
  AND2_X1 U378 ( .A1(net134977), .A2(n85), .ZN(n493) );
  NAND2_X1 U379 ( .A1(\ML_int[7][5] ), .A2(net134975), .ZN(n559) );
  NOR2_X1 U380 ( .A1(n82), .A2(n325), .ZN(\ML_int[7][5] ) );
  NAND2_X1 U381 ( .A1(n433), .A2(n434), .ZN(\ML_int[3][8] ) );
  NAND2_X1 U382 ( .A1(\ML_int[2][8] ), .A2(net134927), .ZN(n433) );
  NAND2_X1 U383 ( .A1(\ML_int[2][4] ), .A2(net134943), .ZN(n434) );
  NAND2_X1 U384 ( .A1(n171), .A2(net134833), .ZN(n607) );
  AND2_X1 U385 ( .A1(\ML_int[4][14] ), .A2(n622), .ZN(\ML_int[7][14] ) );
  CLKBUF_X1 U386 ( .A(net134913), .Z(net134893) );
  NAND2_X1 U387 ( .A1(\MR_int[2][21] ), .A2(net134937), .ZN(n478) );
  NAND2_X1 U388 ( .A1(\ML_int[2][6] ), .A2(net134939), .ZN(n540) );
  NAND2_X1 U390 ( .A1(\ML_int[2][12] ), .A2(net134927), .ZN(n320) );
  NAND2_X1 U391 ( .A1(\ML_int[2][14] ), .A2(net134939), .ZN(n521) );
  NAND2_X1 U392 ( .A1(\ML_int[2][18] ), .A2(net134927), .ZN(net60893) );
  NAND2_X1 U393 ( .A1(\ML_int[2][5] ), .A2(net134925), .ZN(n300) );
  AND2_X1 U394 ( .A1(n85), .A2(net134977), .ZN(n227) );
  AND2_X1 U395 ( .A1(n85), .A2(net134977), .ZN(n379) );
  NAND2_X1 U396 ( .A1(n507), .A2(n506), .ZN(n253) );
  NAND2_X1 U397 ( .A1(\ML_int[2][20] ), .A2(net134927), .ZN(n506) );
  NAND2_X1 U398 ( .A1(n141), .A2(n142), .ZN(\ML_int[3][15] ) );
  NAND2_X1 U399 ( .A1(\ML_int[2][15] ), .A2(net134925), .ZN(n141) );
  NAND2_X1 U400 ( .A1(n538), .A2(n537), .ZN(\ML_int[3][11] ) );
  NAND2_X1 U401 ( .A1(\ML_int[2][7] ), .A2(net134941), .ZN(n538) );
  CLKBUF_X1 U402 ( .A(net134913), .Z(net134891) );
  CLKBUF_X1 U403 ( .A(net134911), .Z(net134899) );
  AND2_X1 U404 ( .A1(net134827), .A2(n85), .ZN(n252) );
  OR2_X1 U405 ( .A1(n271), .A2(net134977), .ZN(n335) );
  NAND2_X1 U406 ( .A1(n345), .A2(n357), .ZN(n355) );
  NAND2_X1 U407 ( .A1(\MR_int[2][23] ), .A2(net134923), .ZN(n545) );
  AND2_X1 U408 ( .A1(\ML_int[2][3] ), .A2(net134925), .ZN(\ML_int[3][3] ) );
  AND2_X1 U409 ( .A1(\ML_int[2][2] ), .A2(net134925), .ZN(\ML_int[3][2] ) );
  NAND2_X1 U410 ( .A1(\ML_int[2][5] ), .A2(net134933), .ZN(n466) );
  NAND2_X1 U411 ( .A1(n517), .A2(n516), .ZN(\ML_int[3][13] ) );
  AND2_X1 U412 ( .A1(\MR_int[3][29] ), .A2(net134843), .ZN(\MR_int[4][29] ) );
  AND2_X1 U413 ( .A1(n623), .A2(n624), .ZN(\MR_int[4][28] ) );
  INV_X1 U414 ( .A(n85), .ZN(n758) );
  CLKBUF_X1 U415 ( .A(net134911), .Z(net134895) );
  NAND2_X1 U416 ( .A1(n220), .A2(n221), .ZN(n225) );
  NOR2_X1 U417 ( .A1(n392), .A2(n162), .ZN(n221) );
  NAND2_X1 U418 ( .A1(net134953), .A2(net61436), .ZN(n162) );
  NAND2_X1 U419 ( .A1(\ML_int[3][27] ), .A2(net134833), .ZN(n430) );
  NAND2_X1 U420 ( .A1(n480), .A2(n481), .ZN(\ML_int[3][27] ) );
  NAND2_X1 U421 ( .A1(n250), .A2(net134923), .ZN(n480) );
  NAND2_X1 U422 ( .A1(\ML_int[2][23] ), .A2(net134951), .ZN(n481) );
  NAND2_X1 U423 ( .A1(net61755), .A2(n349), .ZN(\MR_int[4][6] ) );
  NAND2_X1 U424 ( .A1(\MR_int[3][6] ), .A2(net134849), .ZN(n349) );
  NAND2_X1 U425 ( .A1(\MR_int[3][14] ), .A2(net134831), .ZN(net61755) );
  NAND2_X1 U426 ( .A1(\ML_int[3][24] ), .A2(net134837), .ZN(n431) );
  NAND2_X1 U427 ( .A1(n341), .A2(n342), .ZN(\ML_int[3][24] ) );
  NAND2_X1 U428 ( .A1(\ML_int[2][20] ), .A2(net134933), .ZN(n342) );
  NAND2_X1 U429 ( .A1(n518), .A2(n519), .ZN(\ML_int[3][16] ) );
  NAND2_X1 U430 ( .A1(\ML_int[2][12] ), .A2(net134945), .ZN(n519) );
  NAND2_X1 U431 ( .A1(n410), .A2(net134927), .ZN(n407) );
  NAND2_X1 U432 ( .A1(n484), .A2(n485), .ZN(\MR_int[3][24] ) );
  NAND2_X1 U433 ( .A1(n473), .A2(n474), .ZN(\ML_int[3][7] ) );
  NAND2_X1 U434 ( .A1(\ML_int[2][3] ), .A2(net134943), .ZN(n474) );
  NAND2_X1 U435 ( .A1(\ML_int[2][7] ), .A2(net134925), .ZN(n473) );
  NOR2_X1 U436 ( .A1(n325), .A2(n88), .ZN(\ML_int[7][0] ) );
  NOR2_X1 U437 ( .A1(n325), .A2(n86), .ZN(\ML_int[7][2] ) );
  NOR2_X1 U438 ( .A1(n325), .A2(n87), .ZN(\ML_int[7][1] ) );
  NOR2_X1 U439 ( .A1(n80), .A2(n325), .ZN(\ML_int[7][7] ) );
  AND2_X1 U440 ( .A1(\ML_int[2][0] ), .A2(net134923), .ZN(\ML_int[3][0] ) );
  AND2_X1 U441 ( .A1(\ML_int[2][1] ), .A2(net134925), .ZN(\ML_int[3][1] ) );
  NAND2_X1 U442 ( .A1(n375), .A2(n376), .ZN(\ML_int[7][28] ) );
  NAND2_X1 U443 ( .A1(\ML_int[4][28] ), .A2(n252), .ZN(n376) );
  NAND2_X1 U444 ( .A1(\ML_int[4][12] ), .A2(n377), .ZN(n375) );
  NAND2_X1 U445 ( .A1(n552), .A2(n553), .ZN(\ML_int[3][14] ) );
  NAND2_X1 U446 ( .A1(\ML_int[2][14] ), .A2(net134923), .ZN(n552) );
  NAND2_X1 U447 ( .A1(n489), .A2(n488), .ZN(\ML_int[4][25] ) );
  NAND2_X1 U449 ( .A1(\ML_int[3][25] ), .A2(net134831), .ZN(n488) );
  NAND2_X1 U450 ( .A1(n466), .A2(n465), .ZN(\ML_int[3][9] ) );
  NAND2_X1 U451 ( .A1(\ML_int[3][29] ), .A2(net134831), .ZN(n387) );
  NAND2_X1 U452 ( .A1(\MR_int[2][8] ), .A2(net134935), .ZN(n406) );
  NAND2_X1 U453 ( .A1(\ML_int[2][24] ), .A2(net134935), .ZN(n418) );
  AND2_X1 U454 ( .A1(net134811), .A2(n85), .ZN(n377) );
  AND2_X1 U455 ( .A1(net134811), .A2(n261), .ZN(n234) );
  NAND2_X1 U456 ( .A1(\MR_int[3][18] ), .A2(net134839), .ZN(n575) );
  NAND2_X1 U457 ( .A1(n460), .A2(n461), .ZN(B[6]) );
  NAND2_X1 U458 ( .A1(\MR_int[4][22] ), .A2(n189), .ZN(n428) );
  NOR2_X1 U459 ( .A1(net134971), .A2(net61266), .ZN(n189) );
  OR2_X1 U460 ( .A1(n476), .A2(n180), .ZN(n168) );
  NAND2_X1 U461 ( .A1(\MR_int[4][30] ), .A2(net134969), .ZN(n180) );
  NAND2_X1 U462 ( .A1(n754), .A2(net134809), .ZN(n304) );
  NAND2_X1 U463 ( .A1(n486), .A2(n487), .ZN(\ML_int[3][25] ) );
  NAND2_X1 U464 ( .A1(\ML_int[2][25] ), .A2(net134923), .ZN(n486) );
  NAND2_X1 U465 ( .A1(\ML_int[5][26] ), .A2(n493), .ZN(n525) );
  NAND2_X1 U466 ( .A1(\ML_int[4][26] ), .A2(net134821), .ZN(n298) );
  NAND2_X1 U467 ( .A1(n163), .A2(n164), .ZN(n568) );
  OR2_X1 U468 ( .A1(n746), .A2(n226), .ZN(n164) );
  AND2_X1 U469 ( .A1(net134811), .A2(n306), .ZN(n226) );
  NAND2_X1 U470 ( .A1(n450), .A2(n451), .ZN(B[17]) );
  OR2_X1 U471 ( .A1(n210), .A2(n541), .ZN(n451) );
  NAND2_X1 U472 ( .A1(n525), .A2(n524), .ZN(B[26]) );
  OR2_X1 U473 ( .A1(n388), .A2(net60660), .ZN(n524) );
  NAND2_X1 U474 ( .A1(n156), .A2(n157), .ZN(n572) );
  NOR2_X1 U475 ( .A1(net134969), .A2(net60660), .ZN(n157) );
  NAND2_X1 U476 ( .A1(n427), .A2(n428), .ZN(B[21]) );
  NAND2_X1 U477 ( .A1(\ML_int[3][1] ), .A2(net134853), .ZN(n409) );
  NAND2_X1 U478 ( .A1(n345), .A2(n365), .ZN(n363) );
  NAND2_X1 U479 ( .A1(n181), .A2(net61436), .ZN(n558) );
  NAND2_X1 U480 ( .A1(\ML_int[5][21] ), .A2(net61624), .ZN(n427) );
  AND2_X1 U481 ( .A1(n85), .A2(net134977), .ZN(net61624) );
  NAND2_X1 U482 ( .A1(n124), .A2(n125), .ZN(\ML_int[5][21] ) );
  NAND2_X1 U483 ( .A1(\ML_int[4][21] ), .A2(net134821), .ZN(n124) );
  AND2_X1 U484 ( .A1(n622), .A2(net134977), .ZN(n211) );
  AND2_X1 U485 ( .A1(net134813), .A2(n237), .ZN(n204) );
  AND2_X1 U486 ( .A1(net134813), .A2(n405), .ZN(n241) );
  OR2_X1 U487 ( .A1(n358), .A2(n359), .ZN(n435) );
  NAND2_X1 U488 ( .A1(n223), .A2(net134809), .ZN(n358) );
  NAND2_X1 U489 ( .A1(n738), .A2(n739), .ZN(n454) );
  NAND2_X1 U490 ( .A1(n627), .A2(n628), .ZN(n738) );
  NOR2_X1 U491 ( .A1(net134971), .A2(net61266), .ZN(n739) );
  AND2_X1 U492 ( .A1(\ML_int[4][15] ), .A2(net134977), .ZN(n384) );
  AND2_X1 U494 ( .A1(\ML_int[4][12] ), .A2(net134977), .ZN(n235) );
  NAND2_X1 U495 ( .A1(n272), .A2(n273), .ZN(n499) );
  NAND2_X1 U496 ( .A1(\MR_int[4][25] ), .A2(net134969), .ZN(n412) );
  NAND2_X1 U497 ( .A1(n308), .A2(n307), .ZN(\MR_int[3][12] ) );
  NAND2_X1 U498 ( .A1(n410), .A2(net134951), .ZN(n307) );
  NAND2_X1 U499 ( .A1(net61331), .A2(n439), .ZN(\MR_int[3][10] ) );
  NAND2_X1 U500 ( .A1(\MR_int[2][10] ), .A2(net134953), .ZN(n439) );
  NAND2_X1 U501 ( .A1(n131), .A2(n132), .ZN(\ML_int[5][31] ) );
  NAND2_X1 U502 ( .A1(\ML_int[4][31] ), .A2(net134815), .ZN(n131) );
  NAND2_X1 U503 ( .A1(\ML_int[4][15] ), .A2(net134809), .ZN(n132) );
  AND2_X1 U504 ( .A1(net134971), .A2(n549), .ZN(n201) );
  NAND2_X1 U505 ( .A1(\MR_int[4][28] ), .A2(net134969), .ZN(n592) );
  NAND2_X1 U506 ( .A1(\ML_int[2][25] ), .A2(net134949), .ZN(n390) );
  NAND2_X1 U507 ( .A1(\ML_int[5][30] ), .A2(n421), .ZN(n529) );
  AND2_X1 U508 ( .A1(n85), .A2(net134977), .ZN(n421) );
  AND2_X1 U509 ( .A1(net134811), .A2(n273), .ZN(n214) );
  AND2_X1 U510 ( .A1(net134811), .A2(net61436), .ZN(n170) );
  NAND2_X1 U511 ( .A1(\MR_int[3][16] ), .A2(net134853), .ZN(n627) );
  OR2_X1 U512 ( .A1(net60660), .A2(net134971), .ZN(n210) );
  OR2_X1 U513 ( .A1(n359), .A2(n449), .ZN(n256) );
  AND2_X1 U514 ( .A1(net134859), .A2(net134971), .ZN(n175) );
  OR2_X1 U515 ( .A1(n207), .A2(n208), .ZN(n319) );
  OR2_X1 U516 ( .A1(n748), .A2(net134971), .ZN(n207) );
  INV_X1 U517 ( .A(\MR_int[4][29] ), .ZN(n748) );
  NAND2_X1 U518 ( .A1(\MR_int[4][8] ), .A2(n257), .ZN(n255) );
  AND2_X1 U519 ( .A1(net134811), .A2(n237), .ZN(n257) );
  NAND2_X1 U520 ( .A1(n406), .A2(n407), .ZN(\MR_int[3][8] ) );
  NAND2_X1 U521 ( .A1(n229), .A2(n230), .ZN(n233) );
  NAND2_X1 U522 ( .A1(\MR_int[4][10] ), .A2(n234), .ZN(n232) );
  AND2_X1 U523 ( .A1(n237), .A2(net134971), .ZN(n230) );
  NAND2_X1 U524 ( .A1(\MR_int[4][29] ), .A2(net134969), .ZN(n456) );
  NOR2_X1 U525 ( .A1(\SHMAG[5] ), .A2(net134975), .ZN(net61436) );
  NOR2_X1 U526 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(n237) );
  AND2_X1 U527 ( .A1(n602), .A2(n603), .ZN(n580) );
  NOR2_X1 U528 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(n273) );
  NOR2_X1 U529 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(n405) );
  NOR2_X1 U530 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(n549) );
  NOR2_X1 U531 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(n261) );
  NAND2_X1 U532 ( .A1(n696), .A2(n212), .ZN(B[3]) );
  NOR2_X1 U533 ( .A1(\SHMAG[5] ), .A2(net134975), .ZN(n306) );
  NAND2_X1 U534 ( .A1(\ML_int[1][18] ), .A2(net134891), .ZN(net61783) );
  NAND2_X1 U535 ( .A1(\ML_int[1][10] ), .A2(net134885), .ZN(n483) );
  NAND2_X1 U536 ( .A1(\ML_int[1][5] ), .A2(net134885), .ZN(n441) );
  NAND2_X1 U537 ( .A1(\ML_int[1][6] ), .A2(net134885), .ZN(n492) );
  NOR2_X1 U538 ( .A1(net134971), .A2(\SHMAG[5] ), .ZN(n391) );
  AND2_X1 U539 ( .A1(\MR_int[4][25] ), .A2(n391), .ZN(\MR_int[7][24] ) );
  NAND2_X1 U540 ( .A1(\ML_int[1][19] ), .A2(net134893), .ZN(n459) );
  NAND2_X1 U541 ( .A1(\MR_int[1][7] ), .A2(net134893), .ZN(n398) );
  NAND2_X1 U542 ( .A1(\MR_int[1][14] ), .A2(net134887), .ZN(n282) );
  NAND2_X1 U543 ( .A1(\ML_int[1][16] ), .A2(net134889), .ZN(net60604) );
  NAND2_X1 U544 ( .A1(n200), .A2(n505), .ZN(\ML_int[2][9] ) );
  OR2_X1 U545 ( .A1(net134977), .A2(\SHMAG[5] ), .ZN(n359) );
  NAND2_X1 U546 ( .A1(n728), .A2(net134887), .ZN(n344) );
  NAND2_X1 U547 ( .A1(n508), .A2(n509), .ZN(\ML_int[2][14] ) );
  NAND2_X1 U548 ( .A1(\ML_int[1][12] ), .A2(net134887), .ZN(n509) );
  NAND2_X1 U549 ( .A1(n452), .A2(n453), .ZN(\ML_int[2][25] ) );
  NAND2_X1 U550 ( .A1(\ML_int[1][23] ), .A2(net134887), .ZN(n453) );
  NAND2_X1 U551 ( .A1(n393), .A2(n394), .ZN(\ML_int[2][6] ) );
  NAND2_X1 U552 ( .A1(\MR_int[1][3] ), .A2(net134889), .ZN(n394) );
  NAND2_X1 U553 ( .A1(\ML_int[2][17] ), .A2(net134945), .ZN(n511) );
  NAND2_X1 U554 ( .A1(n457), .A2(n302), .ZN(\ML_int[2][17] ) );
  OR2_X1 U555 ( .A1(net134977), .A2(\SHMAG[5] ), .ZN(net60660) );
  NAND2_X1 U556 ( .A1(\ML_int[1][7] ), .A2(net134883), .ZN(n505) );
  NAND2_X1 U559 ( .A1(n530), .A2(net60869), .ZN(\ML_int[2][4] ) );
  NAND2_X1 U560 ( .A1(\ML_int[1][2] ), .A2(net134897), .ZN(n530) );
  NAND2_X1 U561 ( .A1(n608), .A2(n609), .ZN(\MR_int[2][21] ) );
  NAND2_X1 U562 ( .A1(\MR_int[1][21] ), .A2(net134891), .ZN(n608) );
  NAND2_X1 U563 ( .A1(n195), .A2(n196), .ZN(\ML_int[2][2] ) );
  NAND2_X1 U564 ( .A1(\ML_int[1][0] ), .A2(net134893), .ZN(n196) );
  NAND2_X1 U566 ( .A1(n121), .A2(n122), .ZN(\ML_int[2][23] ) );
  NAND2_X1 U567 ( .A1(\ML_int[1][21] ), .A2(net134885), .ZN(n122) );
  NOR2_X1 U568 ( .A1(\SHMAG[5] ), .A2(n15), .ZN(\MR_int[7][29] ) );
  OR2_X1 U569 ( .A1(net134971), .A2(n743), .ZN(n15) );
  NAND2_X1 U570 ( .A1(n497), .A2(n498), .ZN(\MR_int[2][8] ) );
  NAND2_X1 U571 ( .A1(\MR_int[1][8] ), .A2(net134897), .ZN(n497) );
  NAND2_X1 U572 ( .A1(n591), .A2(n590), .ZN(\MR_int[3][16] ) );
  NAND2_X1 U573 ( .A1(net60588), .A2(net60589), .ZN(\MR_int[3][14] ) );
  OR2_X1 U574 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(net61266) );
  NAND2_X1 U575 ( .A1(n326), .A2(n327), .ZN(\ML_int[2][18] ) );
  NAND2_X1 U576 ( .A1(\MR_int[1][15] ), .A2(net134895), .ZN(n327) );
  NAND2_X1 U577 ( .A1(\ML_int[2][29] ), .A2(net134923), .ZN(n389) );
  NAND2_X1 U578 ( .A1(n413), .A2(n414), .ZN(\ML_int[2][29] ) );
  NAND2_X1 U579 ( .A1(n424), .A2(net134883), .ZN(n413) );
  NAND2_X1 U580 ( .A1(n457), .A2(n302), .ZN(n348) );
  NAND2_X1 U581 ( .A1(n595), .A2(n596), .ZN(\MR_int[2][19] ) );
  MUX2_X1 U582 ( .A(\MR_int[1][11] ), .B(\MR_int[1][9] ), .S(net134903), .Z(
        \MR_int[2][9] ) );
  OR2_X1 U583 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(n208) );
  NAND2_X1 U584 ( .A1(\ML_int[1][17] ), .A2(net134883), .ZN(n353) );
  NAND2_X1 U585 ( .A1(n568), .A2(n569), .ZN(B[14]) );
  NAND2_X1 U586 ( .A1(n420), .A2(n419), .ZN(\ML_int[4][28] ) );
  NAND2_X1 U587 ( .A1(\ML_int[3][28] ), .A2(net134831), .ZN(n419) );
  NAND2_X1 U588 ( .A1(n253), .A2(net134849), .ZN(n420) );
  NAND2_X1 U589 ( .A1(n418), .A2(n417), .ZN(\ML_int[3][28] ) );
  NAND2_X1 U590 ( .A1(n443), .A2(n442), .ZN(B[20]) );
  NOR2_X1 U591 ( .A1(net134975), .A2(\SHMAG[5] ), .ZN(n313) );
  AND2_X1 U592 ( .A1(n182), .A2(n183), .ZN(n534) );
  NAND2_X1 U593 ( .A1(n436), .A2(n435), .ZN(B[18]) );
  NAND2_X1 U594 ( .A1(\ML_int[5][18] ), .A2(n227), .ZN(n436) );
  AND2_X1 U595 ( .A1(\MR_int[4][31] ), .A2(n391), .ZN(\MR_int[7][30] ) );
  AND2_X1 U596 ( .A1(n598), .A2(n597), .ZN(n305) );
  INV_X1 U597 ( .A(\MR_int[1][31] ), .ZN(n747) );
  OR2_X1 U598 ( .A1(\SHMAG[5] ), .A2(net134977), .ZN(n476) );
  NAND2_X1 U599 ( .A1(n311), .A2(n310), .ZN(\ML_int[2][22] ) );
  NAND2_X1 U600 ( .A1(\ML_int[1][20] ), .A2(net134897), .ZN(n310) );
  NAND2_X1 U602 ( .A1(n150), .A2(n151), .ZN(\ML_int[3][31] ) );
  NAND2_X1 U603 ( .A1(n250), .A2(net134935), .ZN(n150) );
  NOR2_X1 U604 ( .A1(n740), .A2(n741), .ZN(\MR_int[7][20] ) );
  AND2_X1 U605 ( .A1(n606), .A2(n607), .ZN(n740) );
  OR2_X1 U606 ( .A1(\SHMAG[5] ), .A2(net134969), .ZN(n741) );
  INV_X1 U607 ( .A(A[31]), .ZN(n749) );
  MUX2_X1 U608 ( .A(A[22]), .B(A[21]), .S(n705), .Z(\MR_int[1][21] ) );
  NAND2_X1 U609 ( .A1(\ML_int[1][15] ), .A2(net134899), .ZN(n302) );
  NAND2_X1 U610 ( .A1(\MR_int[1][22] ), .A2(net134901), .ZN(n561) );
  NAND2_X1 U611 ( .A1(\ML_int[2][28] ), .A2(net134923), .ZN(n417) );
  NAND2_X1 U612 ( .A1(\MR_int[1][2] ), .A2(net134899), .ZN(n154) );
  NAND2_X1 U613 ( .A1(n610), .A2(n611), .ZN(B[1]) );
  NAND2_X1 U614 ( .A1(\ML_int[3][30] ), .A2(net134837), .ZN(n494) );
  AND2_X1 U615 ( .A1(net134925), .A2(net134837), .ZN(n365) );
  AND2_X1 U616 ( .A1(net134837), .A2(n252), .ZN(n158) );
  AND2_X1 U617 ( .A1(net134837), .A2(net134811), .ZN(n246) );
  NAND2_X1 U618 ( .A1(n499), .A2(n500), .ZN(B[8]) );
  BUF_X1 U619 ( .A(\temp_int_SH[0] ), .Z(net135867) );
  CLKBUF_X3 U620 ( .A(net135717), .Z(net135859) );
  NAND2_X1 U622 ( .A1(SH[4]), .A2(net141507), .ZN(n90) );
  NAND2_X1 U623 ( .A1(SH[5]), .A2(net141507), .ZN(n92) );
  NOR2_X1 U624 ( .A1(net141464), .A2(n747), .ZN(\MR_int[2][31] ) );
  OR2_X1 U625 ( .A1(net135859), .A2(n747), .ZN(n392) );
  NAND2_X1 U626 ( .A1(\MR_int[1][31] ), .A2(net135859), .ZN(n598) );
  AND2_X1 U627 ( .A1(\ML_int[1][0] ), .A2(net135859), .ZN(\ML_int[2][0] ) );
  AND2_X1 U628 ( .A1(\ML_int[1][1] ), .A2(net135859), .ZN(\ML_int[2][1] ) );
  NAND2_X1 U629 ( .A1(n228), .A2(net134833), .ZN(n523) );
  NAND2_X1 U630 ( .A1(\ML_int[3][7] ), .A2(net134831), .ZN(n80) );
  NAND2_X1 U631 ( .A1(\ML_int[3][1] ), .A2(net134837), .ZN(n87) );
  NAND2_X1 U632 ( .A1(\ML_int[3][0] ), .A2(net134837), .ZN(n88) );
  NAND2_X1 U633 ( .A1(\ML_int[1][9] ), .A2(net134879), .ZN(n200) );
  NAND2_X1 U634 ( .A1(\ML_int[1][17] ), .A2(net134879), .ZN(n457) );
  NAND2_X1 U635 ( .A1(\ML_int[1][29] ), .A2(net134879), .ZN(n414) );
  NAND2_X1 U636 ( .A1(\ML_int[1][25] ), .A2(net134879), .ZN(n452) );
  NAND2_X1 U637 ( .A1(net61465), .A2(net141444), .ZN(net135734) );
  INV_X1 U638 ( .A(n729), .ZN(n742) );
  NAND2_X1 U639 ( .A1(n312), .A2(n313), .ZN(n460) );
  NAND2_X1 U640 ( .A1(\MR_int[3][31] ), .A2(net134833), .ZN(n603) );
  AND2_X1 U641 ( .A1(net134861), .A2(\MR_int[3][31] ), .ZN(\MR_int[4][31] ) );
  NOR2_X1 U642 ( .A1(net134927), .A2(n392), .ZN(\MR_int[3][31] ) );
  NOR2_X1 U643 ( .A1(net134929), .A2(n215), .ZN(n228) );
  NOR2_X1 U644 ( .A1(net134929), .A2(n305), .ZN(\MR_int[3][29] ) );
  NOR2_X1 U645 ( .A1(net134929), .A2(n305), .ZN(n171) );
  NOR2_X1 U646 ( .A1(net134837), .A2(net134929), .ZN(n624) );
  NAND2_X1 U647 ( .A1(n348), .A2(net134929), .ZN(n496) );
  NAND2_X1 U648 ( .A1(\ML_int[2][24] ), .A2(net134929), .ZN(n341) );
  NAND2_X1 U649 ( .A1(\ML_int[2][31] ), .A2(net134929), .ZN(n151) );
  NAND2_X1 U650 ( .A1(\ML_int[2][13] ), .A2(net134929), .ZN(n516) );
  AND2_X1 U651 ( .A1(net134963), .A2(net134837), .ZN(n357) );
  NAND2_X1 U652 ( .A1(n337), .A2(n338), .ZN(\MR_int[4][13] ) );
  NAND2_X1 U653 ( .A1(net141562), .A2(net134853), .ZN(n337) );
  NAND2_X1 U654 ( .A1(n623), .A2(net134927), .ZN(n484) );
  NAND2_X1 U655 ( .A1(n251), .A2(net134845), .ZN(n400) );
  NAND2_X1 U656 ( .A1(n251), .A2(net134831), .ZN(n415) );
  NAND2_X1 U657 ( .A1(n492), .A2(n334), .ZN(\ML_int[2][8] ) );
  BUF_X1 U658 ( .A(net134967), .Z(net134957) );
  NAND2_X1 U659 ( .A1(n440), .A2(n441), .ZN(\ML_int[2][7] ) );
  NAND2_X1 U660 ( .A1(\ML_int[1][7] ), .A2(net141528), .ZN(n440) );
  NAND2_X1 U661 ( .A1(\MR_int[2][18] ), .A2(net134923), .ZN(net60588) );
  NAND2_X1 U662 ( .A1(n566), .A2(n567), .ZN(\MR_int[3][20] ) );
  NAND2_X1 U663 ( .A1(\MR_int[1][24] ), .A2(net134893), .ZN(n599) );
  NAND2_X1 U664 ( .A1(\MR_int[2][26] ), .A2(net134923), .ZN(net60477) );
  NAND2_X1 U665 ( .A1(n279), .A2(net60477), .ZN(\MR_int[3][22] ) );
  NAND2_X1 U666 ( .A1(net61774), .A2(net134969), .ZN(n332) );
  NOR2_X1 U667 ( .A1(net134971), .A2(n385), .ZN(n274) );
  NAND2_X1 U668 ( .A1(\ML_int[4][10] ), .A2(net134811), .ZN(n299) );
  NAND2_X1 U669 ( .A1(\ML_int[3][10] ), .A2(net134831), .ZN(n138) );
  NAND2_X1 U670 ( .A1(\ML_int[3][10] ), .A2(net134849), .ZN(n370) );
  NAND2_X1 U671 ( .A1(n540), .A2(n539), .ZN(\ML_int[3][10] ) );
  AND2_X1 U672 ( .A1(n622), .A2(\ML_int[4][13] ), .ZN(\ML_int[7][13] ) );
  NAND2_X1 U673 ( .A1(\ML_int[3][5] ), .A2(net134831), .ZN(n82) );
  NAND2_X1 U674 ( .A1(n529), .A2(n528), .ZN(B[30]) );
  NAND2_X1 U675 ( .A1(n144), .A2(n145), .ZN(\ML_int[4][26] ) );
  NAND2_X1 U676 ( .A1(\ML_int[3][26] ), .A2(net134831), .ZN(n144) );
  NAND2_X1 U677 ( .A1(net134861), .A2(n155), .ZN(n743) );
  NAND2_X1 U678 ( .A1(n533), .A2(n534), .ZN(n312) );
  AND2_X1 U679 ( .A1(net60450), .A2(n104), .ZN(n99) );
  NAND2_X1 U680 ( .A1(\ML_int[3][6] ), .A2(net134833), .ZN(n81) );
  NAND2_X1 U681 ( .A1(n587), .A2(n586), .ZN(\ML_int[3][6] ) );
  OAI21_X1 U682 ( .B1(n219), .B2(net134929), .A(n464), .ZN(\ML_int[3][23] ) );
  NAND2_X1 U683 ( .A1(\ML_int[2][23] ), .A2(net134929), .ZN(n464) );
  NOR2_X1 U684 ( .A1(net134831), .A2(n448), .ZN(n520) );
  NAND2_X1 U685 ( .A1(\ML_int[3][21] ), .A2(net134849), .ZN(n386) );
  NAND2_X1 U686 ( .A1(\MR_int[4][4] ), .A2(n214), .ZN(n212) );
  NAND2_X1 U687 ( .A1(n345), .A2(net134927), .ZN(n465) );
  NAND2_X1 U688 ( .A1(\ML_int[2][9] ), .A2(net134945), .ZN(n517) );
  NAND2_X1 U689 ( .A1(n200), .A2(n505), .ZN(n345) );
  NAND2_X1 U690 ( .A1(\MR_int[3][23] ), .A2(net134843), .ZN(n602) );
  NAND2_X1 U691 ( .A1(\MR_int[3][23] ), .A2(n184), .ZN(n182) );
  NAND2_X1 U692 ( .A1(n576), .A2(n577), .ZN(B[2]) );
  NAND2_X1 U693 ( .A1(\MR_int[5][3] ), .A2(n549), .ZN(n576) );
  NAND2_X1 U694 ( .A1(n314), .A2(n315), .ZN(\MR_int[5][3] ) );
  NAND2_X1 U695 ( .A1(\ML_int[2][16] ), .A2(net134937), .ZN(n507) );
  NAND2_X1 U696 ( .A1(\ML_int[2][16] ), .A2(net134925), .ZN(n518) );
  NAND2_X1 U697 ( .A1(n404), .A2(n403), .ZN(\ML_int[2][16] ) );
  NAND2_X1 U698 ( .A1(n478), .A2(n479), .ZN(\MR_int[3][21] ) );
  NAND2_X1 U699 ( .A1(\MR_int[3][21] ), .A2(net134831), .ZN(n338) );
  NAND2_X1 U700 ( .A1(\MR_int[2][20] ), .A2(net134923), .ZN(n591) );
  NAND2_X1 U701 ( .A1(\MR_int[2][20] ), .A2(net134945), .ZN(n566) );
  NAND2_X1 U702 ( .A1(net61724), .A2(n354), .ZN(\MR_int[2][20] ) );
  NAND2_X1 U703 ( .A1(\ML_int[2][10] ), .A2(net134927), .ZN(n539) );
  NAND2_X1 U704 ( .A1(\ML_int[2][10] ), .A2(net134947), .ZN(n553) );
  NAND2_X1 U705 ( .A1(\ML_int[2][11] ), .A2(net134925), .ZN(n537) );
  NAND2_X1 U706 ( .A1(\ML_int[2][11] ), .A2(net134941), .ZN(n142) );
  NAND2_X1 U707 ( .A1(\MR_int[4][2] ), .A2(net134809), .ZN(n588) );
  NAND2_X1 U708 ( .A1(n153), .A2(n154), .ZN(\MR_int[2][2] ) );
  NAND2_X1 U709 ( .A1(\MR_int[1][4] ), .A2(net134879), .ZN(n153) );
  NAND2_X1 U710 ( .A1(n386), .A2(n387), .ZN(\ML_int[4][29] ) );
  NAND2_X1 U711 ( .A1(n390), .A2(n389), .ZN(\ML_int[3][29] ) );
  NAND2_X1 U712 ( .A1(\MR_int[2][29] ), .A2(net134927), .ZN(n147) );
  NAND2_X1 U713 ( .A1(n445), .A2(n444), .ZN(\MR_int[3][23] ) );
  NAND2_X1 U714 ( .A1(\MR_int[2][23] ), .A2(net134933), .ZN(n445) );
  NAND2_X1 U715 ( .A1(\MR_int[3][9] ), .A2(n745), .ZN(n744) );
  AND2_X1 U716 ( .A1(net134833), .A2(net134811), .ZN(n745) );
  NAND2_X1 U717 ( .A1(n318), .A2(n319), .ZN(B[28]) );
  AND2_X1 U718 ( .A1(net141573), .A2(net134837), .ZN(n309) );
  NAND2_X1 U719 ( .A1(\ML_int[3][4] ), .A2(net134843), .ZN(n416) );
  NAND2_X1 U720 ( .A1(\MR_int[1][6] ), .A2(net134899), .ZN(n380) );
  NAND2_X1 U721 ( .A1(n380), .A2(n381), .ZN(\MR_int[2][6] ) );
  NAND2_X1 U722 ( .A1(n730), .A2(n175), .ZN(n449) );
  AND2_X1 U723 ( .A1(\MR_int[3][24] ), .A2(net134843), .ZN(\MR_int[4][24] ) );
  NAND2_X1 U724 ( .A1(n730), .A2(net134837), .ZN(n628) );
  AND2_X1 U725 ( .A1(net134861), .A2(n155), .ZN(\MR_int[4][30] ) );
  NOR2_X1 U726 ( .A1(net134929), .A2(n751), .ZN(n155) );
  INV_X1 U727 ( .A(\MR_int[2][30] ), .ZN(n751) );
  AND2_X1 U728 ( .A1(n352), .A2(n353), .ZN(n219) );
  NAND2_X1 U729 ( .A1(n353), .A2(n352), .ZN(\ML_int[2][19] ) );
  NAND2_X1 U730 ( .A1(\ML_int[1][19] ), .A2(net135859), .ZN(n352) );
  NAND2_X1 U731 ( .A1(\MR_int[2][11] ), .A2(net134951), .ZN(n554) );
  NAND2_X1 U733 ( .A1(\MR_int[3][7] ), .A2(net134851), .ZN(n192) );
  NAND2_X1 U735 ( .A1(n147), .A2(n148), .ZN(\MR_int[3][25] ) );
  NAND2_X1 U736 ( .A1(\MR_int[2][27] ), .A2(net134927), .ZN(n444) );
  NAND2_X1 U737 ( .A1(\MR_int[4][3] ), .A2(net134809), .ZN(n314) );
  NAND2_X1 U738 ( .A1(n554), .A2(n555), .ZN(\MR_int[3][11] ) );
  NAND2_X1 U739 ( .A1(n511), .A2(n510), .ZN(\ML_int[3][21] ) );
  NAND2_X1 U740 ( .A1(n459), .A2(n458), .ZN(\ML_int[2][21] ) );
  NAND2_X1 U741 ( .A1(n725), .A2(net134969), .ZN(n448) );
  NAND2_X1 U742 ( .A1(\MR_int[3][27] ), .A2(net134831), .ZN(n605) );
  NAND2_X1 U743 ( .A1(net61842), .A2(n604), .ZN(n223) );
  NAND2_X1 U744 ( .A1(n395), .A2(n396), .ZN(\ML_int[4][13] ) );
  AND2_X1 U745 ( .A1(n355), .A2(n356), .ZN(n395) );
  NAND2_X1 U746 ( .A1(\ML_int[3][5] ), .A2(net134845), .ZN(n396) );
  NAND2_X1 U747 ( .A1(n300), .A2(n301), .ZN(\ML_int[3][5] ) );
  NAND2_X1 U748 ( .A1(\ML_int[2][1] ), .A2(net134943), .ZN(n301) );
  NAND2_X1 U749 ( .A1(net61783), .A2(net61782), .ZN(\ML_int[2][20] ) );
  NAND2_X1 U750 ( .A1(n556), .A2(n557), .ZN(\MR_int[3][9] ) );
  AND2_X1 U751 ( .A1(net60450), .A2(n104), .ZN(n286) );
  OR2_X1 U752 ( .A1(n267), .A2(net135875), .ZN(n500) );
  NAND2_X1 U753 ( .A1(\MR_int[7][30] ), .A2(net135876), .ZN(n528) );
  NAND2_X1 U754 ( .A1(\MR_int[7][20] ), .A2(net135875), .ZN(n442) );
  NAND2_X1 U755 ( .A1(\MR_int[7][24] ), .A2(net135875), .ZN(n526) );
  NAND2_X1 U756 ( .A1(n425), .A2(n426), .ZN(\ML_int[4][19] ) );
  NAND2_X1 U757 ( .A1(\ML_int[3][19] ), .A2(net134851), .ZN(n429) );
  NAND2_X1 U758 ( .A1(n135), .A2(n136), .ZN(\MR_int[3][1] ) );
  NAND2_X1 U759 ( .A1(\MR_int[1][5] ), .A2(net134895), .ZN(n333) );
  NAND2_X1 U760 ( .A1(\MR_int[4][20] ), .A2(n201), .ZN(n213) );
  NAND2_X1 U761 ( .A1(n522), .A2(n523), .ZN(\MR_int[4][20] ) );
  NAND2_X1 U762 ( .A1(n522), .A2(n523), .ZN(n156) );
  NAND2_X1 U763 ( .A1(\MR_int[3][20] ), .A2(net134839), .ZN(n522) );
  NAND2_X1 U764 ( .A1(n551), .A2(n550), .ZN(\ML_int[4][14] ) );
  NAND2_X1 U765 ( .A1(n494), .A2(net61053), .ZN(\ML_int[4][30] ) );
  NAND2_X1 U766 ( .A1(\MR_int[1][16] ), .A2(net134895), .ZN(n542) );
  NAND2_X1 U767 ( .A1(\MR_int[1][16] ), .A2(net134879), .ZN(n283) );
  NAND2_X1 U769 ( .A1(n542), .A2(net60763), .ZN(\MR_int[2][16] ) );
  NAND2_X1 U770 ( .A1(\MR_int[2][16] ), .A2(net134923), .ZN(n308) );
  NAND2_X1 U771 ( .A1(\MR_int[2][16] ), .A2(net134949), .ZN(n590) );
  NAND2_X1 U772 ( .A1(n535), .A2(n536), .ZN(\MR_int[3][18] ) );
  NAND2_X1 U773 ( .A1(net61353), .A2(net134947), .ZN(n535) );
  NAND2_X1 U774 ( .A1(n398), .A2(n397), .ZN(\ML_int[2][10] ) );
  NOR2_X1 U775 ( .A1(net61363), .A2(net61364), .ZN(n100) );
  NOR2_X1 U776 ( .A1(net61363), .A2(net61364), .ZN(n284) );
  NAND2_X1 U778 ( .A1(n597), .A2(n598), .ZN(\MR_int[2][29] ) );
  NAND2_X1 U779 ( .A1(\MR_int[1][30] ), .A2(net141464), .ZN(n570) );
  AND2_X1 U780 ( .A1(net134901), .A2(\MR_int[1][30] ), .ZN(\MR_int[2][30] ) );
  NAND2_X1 U781 ( .A1(n97), .A2(net135876), .ZN(n91) );
  NAND2_X1 U782 ( .A1(\MR_int[2][1] ), .A2(net134951), .ZN(n136) );
  NAND2_X1 U783 ( .A1(\MR_int[4][18] ), .A2(net134969), .ZN(n589) );
  NAND2_X1 U784 ( .A1(n563), .A2(n562), .ZN(\MR_int[2][26] ) );
  NAND2_X1 U785 ( .A1(n527), .A2(n526), .ZN(B[24]) );
  NAND2_X1 U786 ( .A1(\ML_int[1][14] ), .A2(net134879), .ZN(n508) );
  NAND2_X1 U787 ( .A1(\ML_int[1][14] ), .A2(net134889), .ZN(n404) );
  NAND2_X1 U788 ( .A1(\MR_int[1][25] ), .A2(net134891), .ZN(n543) );
  NAND2_X1 U789 ( .A1(\MR_int[2][9] ), .A2(net134939), .ZN(n556) );
  NAND2_X1 U790 ( .A1(net61046), .A2(n495), .ZN(B[22]) );
  NOR3_X1 U791 ( .A1(net134969), .A2(\SHMAG[5] ), .A3(n580), .ZN(
        \MR_int[7][22] ) );
  NAND2_X1 U792 ( .A1(\MR_int[1][20] ), .A2(net134901), .ZN(net61724) );
  NAND4_X1 U793 ( .A1(n101), .A2(n98), .A3(n99), .A4(n100), .ZN(n97) );
  NAND2_X1 U794 ( .A1(n584), .A2(n585), .ZN(B[10]) );
  AOI22_X1 U795 ( .A1(\MR_int[4][11] ), .A2(n383), .B1(n520), .B2(n261), .ZN(
        n584) );
  NAND2_X1 U796 ( .A1(\ML_int[7][28] ), .A2(net134977), .ZN(n318) );
  NAND2_X1 U797 ( .A1(\ML_int[7][1] ), .A2(net134977), .ZN(n611) );
  NAND2_X1 U798 ( .A1(\ML_int[7][2] ), .A2(net134977), .ZN(n577) );
  NAND2_X1 U799 ( .A1(\ML_int[7][6] ), .A2(net134977), .ZN(n461) );
  NAND2_X1 U800 ( .A1(\ML_int[7][0] ), .A2(net134977), .ZN(n502) );
  NAND2_X1 U801 ( .A1(\ML_int[7][3] ), .A2(net134977), .ZN(n583) );
  NAND2_X1 U802 ( .A1(\ML_int[7][14] ), .A2(net134977), .ZN(n569) );
  NAND2_X1 U803 ( .A1(\ML_int[7][10] ), .A2(net134977), .ZN(n585) );
  NAND2_X1 U804 ( .A1(\ML_int[7][7] ), .A2(net134977), .ZN(n477) );
  NAND2_X1 U805 ( .A1(n560), .A2(n561), .ZN(\MR_int[2][22] ) );
  NAND2_X1 U806 ( .A1(\MR_int[2][22] ), .A2(net134925), .ZN(n536) );
  NAND2_X1 U807 ( .A1(\MR_int[2][22] ), .A2(net134947), .ZN(n279) );
  NAND2_X1 U808 ( .A1(\MR_int[2][15] ), .A2(net134943), .ZN(n346) );
  NAND2_X1 U809 ( .A1(\MR_int[2][15] ), .A2(net134923), .ZN(n555) );
  NAND2_X1 U810 ( .A1(n581), .A2(net60604), .ZN(\MR_int[2][15] ) );
  NAND2_X1 U811 ( .A1(\MR_int[2][5] ), .A2(net134929), .ZN(n135) );
  NAND2_X1 U812 ( .A1(n333), .A2(n334), .ZN(\MR_int[2][5] ) );
  NAND2_X1 U813 ( .A1(n726), .A2(net134843), .ZN(n197) );
  NAND2_X1 U814 ( .A1(n236), .A2(net134831), .ZN(net61842) );
  NAND2_X1 U815 ( .A1(n178), .A2(n255), .ZN(B[7]) );
  NAND2_X1 U816 ( .A1(\MR_int[1][29] ), .A2(net134899), .ZN(n597) );
  NAND2_X1 U817 ( .A1(n347), .A2(n346), .ZN(\MR_int[3][15] ) );
  NAND2_X1 U818 ( .A1(\MR_int[2][24] ), .A2(net134941), .ZN(n485) );
  NAND2_X1 U819 ( .A1(\MR_int[2][24] ), .A2(net134925), .ZN(n567) );
  NAND2_X1 U820 ( .A1(n332), .A2(n331), .ZN(n181) );
  NAND2_X1 U821 ( .A1(\MR_int[4][6] ), .A2(net134809), .ZN(n331) );
  NAND2_X1 U822 ( .A1(\MR_int[2][14] ), .A2(net134947), .ZN(net60589) );
  NAND2_X1 U823 ( .A1(\MR_int[2][14] ), .A2(net134923), .ZN(net61331) );
  NAND2_X1 U824 ( .A1(n283), .A2(n282), .ZN(\MR_int[2][14] ) );
  NAND2_X1 U825 ( .A1(n599), .A2(n600), .ZN(\MR_int[2][24] ) );
  NAND2_X1 U826 ( .A1(\MR_int[1][26] ), .A2(net134895), .ZN(n562) );
  AND2_X1 U827 ( .A1(n578), .A2(n665), .ZN(n224) );
  NAND2_X1 U828 ( .A1(\MR_int[2][25] ), .A2(net134935), .ZN(n148) );
  NAND2_X1 U829 ( .A1(\MR_int[2][25] ), .A2(net134927), .ZN(n479) );
  NAND2_X1 U830 ( .A1(n543), .A2(n544), .ZN(\MR_int[2][25] ) );
  NAND2_X1 U831 ( .A1(\MR_int[3][9] ), .A2(net134843), .ZN(n467) );
  NAND2_X1 U832 ( .A1(\ML_int[3][18] ), .A2(net134833), .ZN(n369) );
  NAND2_X1 U833 ( .A1(n521), .A2(net60893), .ZN(\ML_int[3][18] ) );
  NAND2_X1 U834 ( .A1(\MR_int[1][10] ), .A2(net134875), .ZN(n498) );
  NAND2_X1 U835 ( .A1(\MR_int[1][18] ), .A2(net141528), .ZN(net60763) );
  NAND2_X1 U836 ( .A1(\MR_int[1][8] ), .A2(net141464), .ZN(n381) );
  NAND2_X1 U837 ( .A1(n186), .A2(net134875), .ZN(n354) );
  NAND2_X1 U838 ( .A1(\ML_int[1][4] ), .A2(net135858), .ZN(net60869) );
  NAND2_X1 U839 ( .A1(\ML_int[1][8] ), .A2(net135858), .ZN(n334) );
  NAND2_X1 U840 ( .A1(\ML_int[1][22] ), .A2(net135858), .ZN(n311) );
  NAND2_X1 U841 ( .A1(\ML_int[1][2] ), .A2(net141528), .ZN(n195) );
  NAND2_X1 U842 ( .A1(\ML_int[1][18] ), .A2(net135858), .ZN(n326) );
  NOR2_X1 U843 ( .A1(net60750), .A2(net60751), .ZN(n101) );
  NOR2_X1 U844 ( .A1(net60750), .A2(net60751), .ZN(n285) );
  NAND2_X1 U845 ( .A1(\MR_int[2][21] ), .A2(net134927), .ZN(n565) );
  AND2_X1 U846 ( .A1(n574), .A2(n575), .ZN(n541) );
  NAND2_X1 U847 ( .A1(n660), .A2(n575), .ZN(\MR_int[4][18] ) );
  NAND2_X1 U848 ( .A1(\MR_int[7][22] ), .A2(net135876), .ZN(net61046) );
  NAND2_X1 U849 ( .A1(n564), .A2(n565), .ZN(\MR_int[3][17] ) );
  NAND2_X1 U850 ( .A1(n264), .A2(net134933), .ZN(net61039) );
  NAND2_X1 U851 ( .A1(n496), .A2(net61039), .ZN(\ML_int[3][17] ) );
  NAND2_X1 U852 ( .A1(\ML_int[4][17] ), .A2(net134821), .ZN(n360) );
  NAND2_X1 U853 ( .A1(n351), .A2(n350), .ZN(\ML_int[2][11] ) );
  NAND2_X1 U854 ( .A1(\ML_int[1][9] ), .A2(net134889), .ZN(n351) );
  NAND2_X1 U855 ( .A1(n514), .A2(n515), .ZN(B[23]) );
  NAND2_X1 U856 ( .A1(n571), .A2(n570), .ZN(n623) );
  AND2_X1 U857 ( .A1(n570), .A2(n571), .ZN(n215) );
  NAND2_X1 U858 ( .A1(n336), .A2(n335), .ZN(B[25]) );
  NOR2_X1 U859 ( .A1(net65464), .A2(net65465), .ZN(n98) );
  NOR2_X1 U860 ( .A1(net65464), .A2(net65465), .ZN(n270) );
  NAND2_X1 U861 ( .A1(n411), .A2(n412), .ZN(n272) );
  NAND2_X1 U862 ( .A1(\MR_int[3][17] ), .A2(net134839), .ZN(n579) );
  NAND2_X1 U863 ( .A1(\MR_int[3][15] ), .A2(net134851), .ZN(n422) );
  NAND2_X1 U864 ( .A1(\MR_int[3][15] ), .A2(net134831), .ZN(n193) );
  NAND2_X1 U865 ( .A1(\MR_int[2][19] ), .A2(net134949), .ZN(n546) );
  NAND2_X1 U866 ( .A1(\MR_int[2][19] ), .A2(net134925), .ZN(n347) );
  NAND2_X1 U867 ( .A1(\MR_int[3][25] ), .A2(net134833), .ZN(n243) );
  AND2_X1 U868 ( .A1(\MR_int[3][25] ), .A2(net134839), .ZN(\MR_int[4][25] ) );
  NAND2_X1 U869 ( .A1(\MR_int[3][25] ), .A2(net134833), .ZN(n578) );
  NAND2_X1 U870 ( .A1(\MR_int[1][24] ), .A2(net141528), .ZN(n560) );
  NAND2_X1 U871 ( .A1(n482), .A2(n483), .ZN(\ML_int[2][12] ) );
  NAND2_X1 U872 ( .A1(\ML_int[1][12] ), .A2(net134879), .ZN(n482) );
  NAND2_X1 U873 ( .A1(n321), .A2(n320), .ZN(n251) );
  NAND2_X1 U874 ( .A1(\ML_int[2][8] ), .A2(net134937), .ZN(n321) );
  NAND2_X1 U875 ( .A1(\MR_int[4][19] ), .A2(net134821), .ZN(n315) );
  NAND2_X1 U876 ( .A1(n605), .A2(n604), .ZN(\MR_int[4][19] ) );
  NAND2_X1 U877 ( .A1(\MR_int[3][19] ), .A2(net134839), .ZN(n604) );
  NAND2_X1 U878 ( .A1(n545), .A2(n546), .ZN(\MR_int[3][19] ) );
  NAND2_X1 U879 ( .A1(n558), .A2(n559), .ZN(B[5]) );
  NAND4_X1 U880 ( .A1(n285), .A2(n286), .A3(n284), .A4(n270), .ZN(net60578) );
  NAND2_X1 U881 ( .A1(\ML_int[3][19] ), .A2(net134831), .ZN(n425) );
  NAND2_X1 U882 ( .A1(\ML_int[2][19] ), .A2(net134925), .ZN(n503) );
  AND2_X1 U883 ( .A1(\MR_int[3][26] ), .A2(net134839), .ZN(n229) );
  NAND2_X1 U884 ( .A1(net134855), .A2(\MR_int[3][26] ), .ZN(n385) );
  NAND2_X1 U885 ( .A1(\MR_int[3][26] ), .A2(net134833), .ZN(n574) );
  NAND2_X1 U886 ( .A1(n732), .A2(net134883), .ZN(n571) );
  AND2_X1 U887 ( .A1(net135715), .A2(n90), .ZN(n173) );
  NAND2_X1 U888 ( .A1(\MR_int[1][28] ), .A2(net141528), .ZN(n563) );
  NAND2_X1 U889 ( .A1(net135715), .A2(n90), .ZN(\temp_int_SH[4] ) );
  AND2_X1 U890 ( .A1(n695), .A2(A[0]), .ZN(\ML_int[1][0] ) );
  NOR2_X1 U891 ( .A1(n749), .A2(net141178), .ZN(\MR_int[1][31] ) );
  NAND2_X1 U892 ( .A1(\ML_int[2][21] ), .A2(net134949), .ZN(n487) );
  NAND2_X1 U893 ( .A1(\MR_int[1][26] ), .A2(net135859), .ZN(n600) );
  NAND2_X1 U894 ( .A1(\ML_int[1][16] ), .A2(net134875), .ZN(n403) );
  NAND2_X1 U895 ( .A1(\ML_int[1][23] ), .A2(net134875), .ZN(n121) );
  NAND2_X1 U896 ( .A1(\ML_int[1][6] ), .A2(net135858), .ZN(n393) );
  NAND2_X1 U897 ( .A1(\ML_int[1][11] ), .A2(net135858), .ZN(n350) );
  NAND2_X1 U898 ( .A1(\ML_int[1][20] ), .A2(net135858), .ZN(net61782) );
  NAND2_X1 U899 ( .A1(\ML_int[1][10] ), .A2(net135859), .ZN(n397) );
  NAND2_X1 U900 ( .A1(\MR_int[1][21] ), .A2(net134875), .ZN(n596) );
  NAND2_X1 U901 ( .A1(\MR_int[1][27] ), .A2(net141528), .ZN(n544) );
  NAND2_X1 U902 ( .A1(n601), .A2(net135859), .ZN(n609) );
  NAND2_X1 U903 ( .A1(\ML_int[1][21] ), .A2(net135858), .ZN(n458) );
  INV_X2 U904 ( .A(net134859), .ZN(net134831) );
  AND2_X4 U905 ( .A1(net135715), .A2(n92), .ZN(\SHMAG[5] ) );
  INV_X1 U906 ( .A(net134825), .ZN(net134813) );
  INV_X1 U907 ( .A(\temp_int_SH[4] ), .ZN(net134815) );
  INV_X1 U908 ( .A(\temp_int_SH[4] ), .ZN(net134819) );
  INV_X1 U909 ( .A(\temp_int_SH[4] ), .ZN(net134821) );
  INV_X1 U910 ( .A(\temp_int_SH[4] ), .ZN(net134825) );
  INV_X1 U911 ( .A(\temp_int_SH[4] ), .ZN(net134827) );
endmodule


module SHIFTER_M32_N5_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [31:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n201, n202, n203, n204, n205, n206, n208, n209, n210, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n240, n241, n242, n243, n244, n245, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n260, n261,
         n263, n265, n266, n268, n272, n273, n279, n280, n283, n286, n287,
         n290, n291, n294, n295, n298, n299, n302, n303, n305, n306, n309,
         n310, n314, n315, n316, n317, n318, n321, n322, n325, n326, n327,
         n329, n330, n331, n332, n334, n335, n336, n337, n338, n341, n342,
         n343, n344, n347, n348, n350, n351, n352, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n371, n372, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n385, n387, n388, n424, n477, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698;

  NAND3_X1 U93 ( .A1(n585), .A2(n696), .A3(n102), .ZN(n100) );
  MUX2_X1 U96 ( .A(n109), .B(n110), .S(n111), .Z(n108) );
  MUX2_X1 U98 ( .A(n115), .B(n116), .S(n111), .Z(n114) );
  MUX2_X1 U100 ( .A(n119), .B(n120), .S(n111), .Z(n118) );
  MUX2_X1 U102 ( .A(n123), .B(n124), .S(n111), .Z(n122) );
  MUX2_X1 U104 ( .A(n127), .B(n128), .S(n111), .Z(n126) );
  MUX2_X1 U106 ( .A(n577), .B(n131), .S(n111), .Z(n129) );
  NAND3_X1 U109 ( .A1(n136), .A2(n137), .A3(n132), .ZN(n135) );
  NAND3_X1 U132 ( .A1(n585), .A2(n696), .A3(n170), .ZN(n177) );
  MUX2_X1 U141 ( .A(n182), .B(n183), .S(n111), .Z(n181) );
  NAND3_X1 U197 ( .A1(n136), .A2(n137), .A3(n206), .ZN(n208) );
  MUX2_X1 U244 ( .A(n189), .B(n190), .S(n111), .Z(n227) );
  NAND3_X1 U23 ( .A1(n290), .A2(n291), .A3(n204), .ZN(n263) );
  NAND3_X1 U46 ( .A1(n351), .A2(n350), .A3(n197), .ZN(n142) );
  NAND3_X1 U59 ( .A1(n279), .A2(n280), .A3(n212), .ZN(n162) );
  NAND3_X1 U71 ( .A1(n286), .A2(n287), .A3(n198), .ZN(n144) );
  NAND3_X1 U76 ( .A1(n290), .A2(n291), .A3(n204), .ZN(n149) );
  NAND3_X1 U81 ( .A1(n294), .A2(n295), .A3(n233), .ZN(n152) );
  NAND3_X1 U86 ( .A1(n298), .A2(n299), .A3(n225), .ZN(n176) );
  NAND3_X1 U94 ( .A1(n302), .A2(n303), .A3(n236), .ZN(n158) );
  NAND3_X1 U107 ( .A1(n305), .A2(n306), .A3(n199), .ZN(n148) );
  NAND3_X1 U122 ( .A1(n314), .A2(n315), .A3(n232), .ZN(n157) );
  NAND3_X1 U130 ( .A1(n224), .A2(n338), .A3(n337), .ZN(n321) );
  NAND3_X1 U138 ( .A1(n325), .A2(n326), .A3(n203), .ZN(n145) );
  NAND3_X1 U154 ( .A1(n337), .A2(n338), .A3(n224), .ZN(n172) );
  NAND3_X1 U170 ( .A1(n347), .A2(n348), .A3(n223), .ZN(n169) );
  NAND3_X1 U182 ( .A1(n358), .A2(n359), .A3(n217), .ZN(n164) );
  NAND3_X1 U190 ( .A1(n365), .A2(n366), .A3(n216), .ZN(n167) );
  NAND3_X1 U193 ( .A1(n367), .A2(n368), .A3(n235), .ZN(n150) );
  NAND3_X1 U200 ( .A1(n371), .A2(n372), .A3(n202), .ZN(n141) );
  NAND3_X1 U208 ( .A1(n215), .A2(n380), .A3(n379), .ZN(n163) );
  NAND3_X1 U373 ( .A1(SH[15]), .A2(SH[14]), .A3(SH[16]), .ZN(n506) );
  NAND2_X2 U281 ( .A1(SH[4]), .A2(n228), .ZN(n111) );
  BUF_X1 U3 ( .A(n273), .Z(n596) );
  CLKBUF_X1 U4 ( .A(n240), .Z(n566) );
  CLKBUF_X3 U5 ( .A(n272), .Z(n639) );
  CLKBUF_X2 U6 ( .A(n272), .Z(n638) );
  OAI221_X1 U7 ( .B1(n616), .B2(n680), .C1(n620), .C2(n676), .A(n219), .ZN(
        n175) );
  BUF_X2 U8 ( .A(n261), .Z(n641) );
  OR2_X1 U9 ( .A1(n694), .A2(n218), .ZN(n113) );
  NOR3_X1 U10 ( .A1(n588), .A2(n589), .A3(n590), .ZN(n131) );
  AND2_X1 U11 ( .A1(n164), .A2(n643), .ZN(n330) );
  AND3_X1 U12 ( .A1(n481), .A2(n482), .A3(n180), .ZN(n105) );
  AOI22_X1 U13 ( .A1(A[30]), .A2(n637), .B1(n639), .B2(A[31]), .ZN(n117) );
  BUF_X2 U14 ( .A(n261), .Z(n643) );
  NOR3_X1 U15 ( .A1(n608), .A2(n609), .A3(n655), .ZN(n134) );
  CLKBUF_X1 U16 ( .A(n240), .Z(n567) );
  AND2_X2 U17 ( .A1(n344), .A2(SH[1]), .ZN(n383) );
  BUF_X1 U18 ( .A(n155), .Z(n568) );
  CLKBUF_X1 U19 ( .A(n145), .Z(n569) );
  AND4_X1 U20 ( .A1(n247), .A2(SH[22]), .A3(SH[20]), .A4(SH[21]), .ZN(n244) );
  OR2_X1 U21 ( .A1(n268), .A2(n690), .ZN(n570) );
  NAND3_X1 U22 ( .A1(n317), .A2(n318), .A3(n221), .ZN(n571) );
  OAI221_X1 U24 ( .B1(n594), .B2(n689), .C1(n619), .C2(n684), .A(n231), .ZN(
        n572) );
  AOI22_X1 U25 ( .A1(A[24]), .A2(n638), .B1(A[25]), .B2(n631), .ZN(n573) );
  BUF_X1 U26 ( .A(n273), .Z(n595) );
  NAND2_X1 U27 ( .A1(n155), .A2(n627), .ZN(n574) );
  NAND2_X1 U28 ( .A1(n158), .A2(n641), .ZN(n575) );
  NAND2_X1 U29 ( .A1(n574), .A2(n575), .ZN(n576) );
  NOR2_X1 U30 ( .A1(n424), .A2(n576), .ZN(n577) );
  BUF_X2 U31 ( .A(n385), .Z(n578) );
  NAND2_X1 U32 ( .A1(n624), .A2(A[15]), .ZN(n336) );
  AOI222_X4 U33 ( .A1(n578), .A2(A[1]), .B1(n638), .B2(A[0]), .C1(n598), .C2(
        A[2]), .ZN(n106) );
  MUX2_X1 U34 ( .A(n160), .B(n159), .S(n196), .Z(n136) );
  OAI221_X1 U35 ( .B1(n693), .B2(n94), .C1(n691), .C2(n93), .A(n570), .ZN(B[7]) );
  AND3_X1 U36 ( .A1(n336), .A2(n335), .A3(n230), .ZN(n266) );
  OAI22_X1 U37 ( .A1(n615), .A2(n579), .B1(n106), .B2(n580), .ZN(n581) );
  INV_X1 U38 ( .A(n600), .ZN(n579) );
  INV_X1 U39 ( .A(n261), .ZN(n580) );
  INV_X1 U40 ( .A(n581), .ZN(n94) );
  NAND2_X1 U41 ( .A1(n584), .A2(n566), .ZN(n273) );
  OAI22_X1 U42 ( .A1(n266), .A2(n615), .B1(n582), .B2(n614), .ZN(n668) );
  INV_X1 U43 ( .A(n153), .ZN(n582) );
  NAND3_X1 U44 ( .A1(n336), .A2(n335), .A3(n230), .ZN(n154) );
  NAND3_X1 U45 ( .A1(n209), .A2(n343), .A3(n342), .ZN(n159) );
  NAND3_X1 U47 ( .A1(n364), .A2(n363), .A3(n362), .ZN(n648) );
  BUF_X1 U48 ( .A(n161), .Z(n583) );
  AND2_X1 U49 ( .A1(n165), .A2(n612), .ZN(n268) );
  INV_X1 U50 ( .A(n383), .ZN(n584) );
  CLKBUF_X1 U51 ( .A(n101), .Z(n585) );
  NAND3_X1 U52 ( .A1(n331), .A2(n332), .A3(n210), .ZN(n586) );
  NAND3_X1 U53 ( .A1(n294), .A2(n295), .A3(n233), .ZN(n587) );
  AND2_X1 U54 ( .A1(n152), .A2(n642), .ZN(n588) );
  AND2_X1 U55 ( .A1(n153), .A2(n626), .ZN(n589) );
  AND2_X1 U56 ( .A1(n157), .A2(n628), .ZN(n590) );
  OR2_X1 U57 ( .A1(n567), .A2(n698), .ZN(n591) );
  OR2_X1 U58 ( .A1(n567), .A2(n698), .ZN(n334) );
  NAND3_X1 U60 ( .A1(n358), .A2(n359), .A3(n217), .ZN(n592) );
  BUF_X1 U61 ( .A(n240), .Z(n604) );
  CLKBUF_X1 U62 ( .A(SH[17]), .Z(n593) );
  INV_X1 U63 ( .A(n165), .ZN(n660) );
  CLKBUF_X1 U64 ( .A(n273), .Z(n594) );
  CLKBUF_X3 U65 ( .A(n272), .Z(n640) );
  INV_X1 U66 ( .A(n334), .ZN(n597) );
  INV_X1 U67 ( .A(n591), .ZN(n598) );
  INV_X1 U68 ( .A(n591), .ZN(n599) );
  INV_X1 U69 ( .A(n334), .ZN(n624) );
  NAND3_X1 U70 ( .A1(n279), .A2(n280), .A3(n212), .ZN(n600) );
  OAI221_X1 U72 ( .B1(n616), .B2(n659), .C1(n656), .C2(n620), .A(n214), .ZN(
        n601) );
  NAND3_X1 U73 ( .A1(n215), .A2(n380), .A3(n379), .ZN(n602) );
  CLKBUF_X1 U74 ( .A(n142), .Z(n603) );
  AND2_X1 U75 ( .A1(n148), .A2(n628), .ZN(n605) );
  AND2_X1 U77 ( .A1(n144), .A2(n642), .ZN(n606) );
  AND2_X1 U78 ( .A1(n137), .A2(n101), .ZN(n607) );
  NOR3_X1 U79 ( .A1(n605), .A2(n606), .A3(n607), .ZN(n128) );
  BUF_X1 U80 ( .A(n385), .Z(n630) );
  AND2_X1 U82 ( .A1(n592), .A2(n627), .ZN(n608) );
  AND2_X1 U83 ( .A1(n167), .A2(n641), .ZN(n609) );
  AND2_X1 U84 ( .A1(n240), .A2(n383), .ZN(n385) );
  AND4_X1 U85 ( .A1(n249), .A2(SH[9]), .A3(SH[7]), .A4(SH[8]), .ZN(n610) );
  CLKBUF_X1 U87 ( .A(SH[28]), .Z(n611) );
  AND4_X1 U88 ( .A1(n249), .A2(SH[9]), .A3(SH[7]), .A4(SH[8]), .ZN(n242) );
  MUX2_X2 U89 ( .A(n142), .B(n143), .S(n196), .Z(n101) );
  NOR2_X1 U90 ( .A1(n330), .A2(n329), .ZN(n612) );
  BUF_X2 U91 ( .A(n385), .Z(n613) );
  INV_X4 U92 ( .A(n102), .ZN(n693) );
  INV_X2 U95 ( .A(n132), .ZN(n690) );
  INV_X2 U97 ( .A(n614), .ZN(n634) );
  INV_X1 U99 ( .A(n614), .ZN(n633) );
  INV_X1 U101 ( .A(n170), .ZN(n692) );
  NAND2_X1 U103 ( .A1(n170), .A2(n628), .ZN(n179) );
  NAND2_X1 U105 ( .A1(n132), .A2(n633), .ZN(n112) );
  INV_X1 U108 ( .A(n615), .ZN(n628) );
  OAI222_X1 U110 ( .A1(n89), .A2(n693), .B1(n91), .B2(n692), .C1(n90), .C2(
        n690), .ZN(B[24]) );
  NOR2_X1 U111 ( .A1(n107), .A2(n695), .ZN(n132) );
  INV_X1 U112 ( .A(n206), .ZN(n691) );
  BUF_X2 U113 ( .A(n387), .Z(n625) );
  NOR2_X1 U114 ( .A1(n113), .A2(n695), .ZN(n170) );
  BUF_X2 U115 ( .A(n385), .Z(n631) );
  BUF_X2 U116 ( .A(n387), .Z(n626) );
  OAI222_X1 U117 ( .A1(n103), .A2(n691), .B1(n683), .B2(n104), .C1(n105), .C2(
        n690), .ZN(B[4]) );
  OAI222_X1 U118 ( .A1(n86), .A2(n690), .B1(n87), .B2(n691), .C1(n88), .C2(
        n693), .ZN(B[9]) );
  OAI221_X1 U119 ( .B1(n98), .B2(n691), .C1(n99), .C2(n690), .A(n100), .ZN(
        B[5]) );
  OAI222_X1 U120 ( .A1(n577), .A2(n690), .B1(n644), .B2(n191), .C1(n131), .C2(
        n693), .ZN(B[12]) );
  OAI222_X1 U121 ( .A1(n138), .A2(n690), .B1(n140), .B2(n691), .C1(n139), .C2(
        n693), .ZN(B[10]) );
  BUF_X2 U123 ( .A(n261), .Z(n642) );
  BUF_X2 U124 ( .A(n387), .Z(n627) );
  BUF_X2 U125 ( .A(n385), .Z(n632) );
  OR2_X2 U126 ( .A1(n697), .A2(n696), .ZN(n614) );
  NAND2_X1 U127 ( .A1(n102), .A2(n628), .ZN(n104) );
  NOR3_X1 U128 ( .A1(n381), .A2(n382), .A3(n651), .ZN(n119) );
  NAND2_X1 U129 ( .A1(n206), .A2(n633), .ZN(n191) );
  OAI222_X1 U131 ( .A1(n92), .A2(n693), .B1(n94), .B2(n692), .C1(n93), .C2(
        n690), .ZN(B[23]) );
  OAI222_X1 U133 ( .A1(n86), .A2(n693), .B1(n88), .B2(n692), .C1(n87), .C2(
        n690), .ZN(B[25]) );
  INV_X1 U134 ( .A(n143), .ZN(n688) );
  OAI222_X1 U135 ( .A1(n95), .A2(n690), .B1(n96), .B2(n691), .C1(n97), .C2(
        n693), .ZN(B[6]) );
  OAI222_X1 U136 ( .A1(n183), .A2(n693), .B1(n688), .B2(n179), .C1(n182), .C2(
        n690), .ZN(B[17]) );
  OAI222_X1 U137 ( .A1(n138), .A2(n693), .B1(n139), .B2(n692), .C1(n140), .C2(
        n690), .ZN(B[26]) );
  OAI221_X1 U139 ( .B1(n99), .B2(n693), .C1(n98), .C2(n690), .A(n177), .ZN(
        B[21]) );
  AND3_X1 U140 ( .A1(n192), .A2(n674), .A3(n679), .ZN(n352) );
  INV_X1 U142 ( .A(n377), .ZN(n679) );
  INV_X1 U143 ( .A(n378), .ZN(n674) );
  INV_X1 U144 ( .A(n160), .ZN(n645) );
  NOR2_X1 U145 ( .A1(n107), .A2(n227), .ZN(B[0]) );
  AOI222_X1 U146 ( .A1(n647), .A2(n643), .B1(n571), .B2(n626), .C1(n169), .C2(
        n633), .ZN(n96) );
  AOI222_X1 U147 ( .A1(n171), .A2(n643), .B1(n687), .B2(n626), .C1(n175), .C2(
        n628), .ZN(n139) );
  AOI222_X1 U148 ( .A1(n159), .A2(n626), .B1(n643), .B2(n160), .C1(n161), .C2(
        n633), .ZN(n93) );
  AOI222_X1 U149 ( .A1(n151), .A2(n642), .B1(n150), .B2(n626), .C1(n158), .C2(
        n633), .ZN(n103) );
  AOI222_X1 U150 ( .A1(n648), .A2(n642), .B1(n141), .B2(n626), .C1(n263), .C2(
        n633), .ZN(n98) );
  OAI22_X1 U151 ( .A1(n615), .A2(n265), .B1(n614), .B2(n266), .ZN(n424) );
  AND3_X1 U152 ( .A1(n367), .A2(n368), .A3(n235), .ZN(n265) );
  AOI221_X1 U153 ( .B1(n152), .B2(n627), .C1(n157), .C2(n641), .A(n668), .ZN(
        n190) );
  NOR2_X1 U155 ( .A1(n113), .A2(n111), .ZN(n102) );
  AOI22_X1 U156 ( .A1(n571), .A2(n633), .B1(n647), .B2(n626), .ZN(n140) );
  AOI22_X1 U157 ( .A1(n141), .A2(n633), .B1(n648), .B2(n626), .ZN(n87) );
  AOI22_X1 U158 ( .A1(n150), .A2(n633), .B1(n151), .B2(n626), .ZN(n90) );
  AOI22_X1 U159 ( .A1(n171), .A2(n628), .B1(n687), .B2(n642), .ZN(n97) );
  NOR2_X1 U160 ( .A1(n107), .A2(n111), .ZN(n206) );
  NAND2_X1 U161 ( .A1(n218), .A2(n694), .ZN(n107) );
  NOR2_X1 U162 ( .A1(n635), .A2(n646), .ZN(n160) );
  AOI22_X1 U163 ( .A1(n634), .A2(n686), .B1(n629), .B2(n602), .ZN(n192) );
  OAI222_X1 U164 ( .A1(n89), .A2(n690), .B1(n90), .B2(n691), .C1(n91), .C2(
        n693), .ZN(B[8]) );
  OAI22_X1 U165 ( .A1(n125), .A2(n112), .B1(n126), .B2(n113), .ZN(B[29]) );
  INV_X1 U166 ( .A(n193), .ZN(n649) );
  AOI22_X1 U167 ( .A1(n634), .A2(n592), .B1(n629), .B2(n159), .ZN(n193) );
  NOR2_X1 U168 ( .A1(n689), .A2(n621), .ZN(n143) );
  INV_X1 U169 ( .A(n106), .ZN(n686) );
  AND3_X1 U171 ( .A1(n483), .A2(n484), .A3(n178), .ZN(n99) );
  NAND2_X1 U172 ( .A1(n569), .A2(n642), .ZN(n484) );
  NAND2_X1 U173 ( .A1(n148), .A2(n625), .ZN(n483) );
  AOI22_X1 U174 ( .A1(n634), .A2(n144), .B1(n628), .B2(n146), .ZN(n178) );
  AOI22_X1 U175 ( .A1(n634), .A2(n602), .B1(n601), .B2(n628), .ZN(n213) );
  AND3_X1 U176 ( .A1(n495), .A2(n496), .A3(n201), .ZN(n127) );
  NAND2_X1 U177 ( .A1(n149), .A2(n641), .ZN(n496) );
  NAND2_X1 U178 ( .A1(n146), .A2(n625), .ZN(n495) );
  AOI22_X1 U179 ( .A1(n634), .A2(n145), .B1(n629), .B2(n141), .ZN(n201) );
  NAND2_X1 U180 ( .A1(n157), .A2(n625), .ZN(n481) );
  AOI22_X1 U181 ( .A1(n634), .A2(n587), .B1(n155), .B2(n628), .ZN(n180) );
  AND3_X1 U183 ( .A1(n186), .A2(n260), .A3(n477), .ZN(n124) );
  NAND2_X1 U184 ( .A1(n172), .A2(n642), .ZN(n260) );
  NAND2_X1 U185 ( .A1(n175), .A2(n625), .ZN(n477) );
  AOI22_X1 U186 ( .A1(n634), .A2(n171), .B1(n629), .B2(n173), .ZN(n186) );
  AND3_X1 U187 ( .A1(n487), .A2(n488), .A3(n174), .ZN(n95) );
  NAND2_X1 U188 ( .A1(n173), .A2(n641), .ZN(n488) );
  NAND2_X1 U189 ( .A1(n321), .A2(n625), .ZN(n487) );
  AOI22_X1 U191 ( .A1(n175), .A2(n633), .B1(n628), .B2(n176), .ZN(n174) );
  OAI22_X1 U192 ( .A1(n108), .A2(n107), .B1(n104), .B2(n106), .ZN(B[3]) );
  OR2_X1 U194 ( .A1(n196), .A2(n137), .ZN(n615) );
  NOR3_X1 U195 ( .A1(n376), .A2(n375), .A3(n374), .ZN(n109) );
  AND2_X1 U196 ( .A1(n192), .A2(n310), .ZN(n116) );
  NOR3_X1 U198 ( .A1(n356), .A2(n357), .A3(n649), .ZN(n115) );
  NOR2_X1 U199 ( .A1(n378), .A2(n377), .ZN(n310) );
  INV_X1 U201 ( .A(n121), .ZN(n687) );
  INV_X1 U202 ( .A(n117), .ZN(n647) );
  INV_X1 U203 ( .A(n151), .ZN(n644) );
  INV_X1 U204 ( .A(n111), .ZN(n695) );
  AND3_X1 U205 ( .A1(n485), .A2(n486), .A3(n147), .ZN(n86) );
  NAND2_X1 U206 ( .A1(n569), .A2(n625), .ZN(n485) );
  NAND2_X1 U207 ( .A1(n146), .A2(n642), .ZN(n486) );
  AOI22_X1 U209 ( .A1(n634), .A2(n148), .B1(n629), .B2(n149), .ZN(n147) );
  AND3_X1 U210 ( .A1(n489), .A2(n490), .A3(n156), .ZN(n89) );
  NAND2_X1 U211 ( .A1(n568), .A2(n641), .ZN(n490) );
  AOI22_X1 U212 ( .A1(n634), .A2(n157), .B1(n628), .B2(n158), .ZN(n156) );
  AND3_X1 U213 ( .A1(n491), .A2(n492), .A3(n222), .ZN(n138) );
  NAND2_X1 U214 ( .A1(n173), .A2(n625), .ZN(n491) );
  NAND2_X1 U215 ( .A1(n176), .A2(n641), .ZN(n492) );
  AOI22_X1 U216 ( .A1(n634), .A2(n321), .B1(n629), .B2(n169), .ZN(n222) );
  AND2_X1 U217 ( .A1(n601), .A2(n627), .ZN(n375) );
  AND2_X1 U218 ( .A1(n169), .A2(n643), .ZN(n382) );
  AND2_X1 U219 ( .A1(n176), .A2(n627), .ZN(n381) );
  OAI222_X1 U220 ( .A1(n95), .A2(n693), .B1(n97), .B2(n692), .C1(n96), .C2(
        n690), .ZN(B[22]) );
  OAI22_X1 U221 ( .A1(n121), .A2(n104), .B1(n107), .B2(n122), .ZN(B[2]) );
  OAI22_X1 U222 ( .A1(n644), .A2(n112), .B1(n113), .B2(n129), .ZN(B[28]) );
  AND2_X1 U223 ( .A1(n162), .A2(n627), .ZN(n377) );
  AND2_X1 U224 ( .A1(n166), .A2(n643), .ZN(n378) );
  INV_X1 U225 ( .A(n195), .ZN(n651) );
  AND3_X1 U226 ( .A1(n493), .A2(n494), .A3(n185), .ZN(n123) );
  NAND2_X1 U227 ( .A1(n168), .A2(n641), .ZN(n494) );
  NAND2_X1 U228 ( .A1(n169), .A2(n625), .ZN(n493) );
  AOI22_X1 U229 ( .A1(n634), .A2(n176), .B1(n629), .B2(n647), .ZN(n185) );
  AND3_X1 U230 ( .A1(n497), .A2(n498), .A3(n188), .ZN(n183) );
  NAND2_X1 U231 ( .A1(n144), .A2(n625), .ZN(n497) );
  NAND2_X1 U232 ( .A1(n148), .A2(n641), .ZN(n498) );
  AND3_X1 U233 ( .A1(n499), .A2(n500), .A3(n184), .ZN(n110) );
  NAND2_X1 U234 ( .A1(n586), .A2(n625), .ZN(n499) );
  NAND2_X1 U235 ( .A1(n602), .A2(n641), .ZN(n500) );
  AND3_X1 U236 ( .A1(n503), .A2(n504), .A3(n194), .ZN(n120) );
  NAND2_X1 U237 ( .A1(n171), .A2(n625), .ZN(n503) );
  NAND2_X1 U238 ( .A1(n175), .A2(n641), .ZN(n504) );
  AOI22_X1 U239 ( .A1(n634), .A2(n687), .B1(n629), .B2(n172), .ZN(n194) );
  AND2_X1 U240 ( .A1(n583), .A2(n643), .ZN(n357) );
  AND2_X1 U241 ( .A1(n327), .A2(n187), .ZN(n182) );
  AOI22_X1 U242 ( .A1(n634), .A2(n146), .B1(n629), .B2(n648), .ZN(n187) );
  NOR2_X1 U243 ( .A1(n360), .A2(n361), .ZN(n327) );
  AND2_X1 U245 ( .A1(n263), .A2(n627), .ZN(n360) );
  AND3_X1 U246 ( .A1(n501), .A2(n502), .A3(n234), .ZN(n189) );
  NAND2_X1 U247 ( .A1(n151), .A2(n628), .ZN(n502) );
  NAND2_X1 U248 ( .A1(n568), .A2(n633), .ZN(n501) );
  AOI22_X1 U249 ( .A1(n626), .A2(n158), .B1(n643), .B2(n150), .ZN(n234) );
  AND2_X1 U250 ( .A1(n163), .A2(n627), .ZN(n329) );
  OAI222_X1 U251 ( .A1(n316), .A2(n690), .B1(n117), .B2(n191), .C1(n693), .C2(
        n120), .ZN(B[14]) );
  NOR3_X1 U252 ( .A1(n381), .A2(n382), .A3(n651), .ZN(n316) );
  OAI222_X1 U253 ( .A1(n105), .A2(n693), .B1(n683), .B2(n179), .C1(n103), .C2(
        n690), .ZN(B[20]) );
  OAI222_X1 U254 ( .A1(n124), .A2(n693), .B1(n121), .B2(n179), .C1(n123), .C2(
        n690), .ZN(B[18]) );
  INV_X1 U255 ( .A(n196), .ZN(n697) );
  AND2_X1 U256 ( .A1(n141), .A2(n643), .ZN(n361) );
  OAI222_X1 U257 ( .A1(n110), .A2(n693), .B1(n106), .B2(n179), .C1(n341), .C2(
        n690), .ZN(B[19]) );
  NOR3_X1 U258 ( .A1(n376), .A2(n375), .A3(n374), .ZN(n341) );
  OR2_X1 U259 ( .A1(n654), .A2(n620), .ZN(n368) );
  OR2_X1 U260 ( .A1(n623), .A2(n671), .ZN(n338) );
  OR2_X1 U261 ( .A1(n622), .A2(n658), .ZN(n291) );
  OR2_X1 U262 ( .A1(n635), .A2(n675), .ZN(n337) );
  OAI221_X1 U263 ( .B1(n616), .B2(n685), .C1(n618), .C2(n681), .A(n220), .ZN(
        n171) );
  OAI221_X1 U264 ( .B1(n635), .B2(n666), .C1(n619), .C2(n663), .A(n205), .ZN(
        n146) );
  AOI22_X1 U265 ( .A1(A[18]), .A2(n640), .B1(A[19]), .B2(n578), .ZN(n205) );
  OAI221_X1 U266 ( .B1(n616), .B2(n667), .C1(n620), .C2(n664), .A(n238), .ZN(
        n155) );
  AOI22_X1 U267 ( .A1(A[17]), .A2(n640), .B1(A[18]), .B2(n631), .ZN(n238) );
  AOI22_X1 U268 ( .A1(A[7]), .A2(n639), .B1(A[8]), .B2(n632), .ZN(n219) );
  OAI221_X1 U269 ( .B1(n594), .B2(n653), .C1(n646), .C2(n622), .A(n237), .ZN(
        n151) );
  AOI22_X1 U270 ( .A1(A[29]), .A2(n639), .B1(n630), .B2(A[30]), .ZN(n237) );
  OR2_X1 U271 ( .A1(n622), .A2(n672), .ZN(n306) );
  AOI22_X1 U272 ( .A1(A[21]), .A2(n640), .B1(A[22]), .B2(n632), .ZN(n236) );
  OR2_X1 U273 ( .A1(n618), .A2(n659), .ZN(n303) );
  AOI22_X1 U274 ( .A1(A[6]), .A2(n640), .B1(A[7]), .B2(n578), .ZN(n198) );
  OR2_X1 U275 ( .A1(n619), .A2(n677), .ZN(n287) );
  AOI22_X1 U276 ( .A1(A[12]), .A2(n638), .B1(A[13]), .B2(n578), .ZN(n215) );
  OR2_X1 U277 ( .A1(n621), .A2(n670), .ZN(n380) );
  OR2_X1 U278 ( .A1(n596), .A2(n665), .ZN(n298) );
  AOI22_X1 U279 ( .A1(A[19]), .A2(n640), .B1(A[20]), .B2(n631), .ZN(n225) );
  OR2_X1 U280 ( .A1(n619), .A2(n662), .ZN(n299) );
  AOI22_X1 U282 ( .A1(A[26]), .A2(n639), .B1(A[27]), .B2(n631), .ZN(n202) );
  OR2_X1 U283 ( .A1(n623), .A2(n653), .ZN(n372) );
  OR2_X1 U284 ( .A1(n622), .A2(n673), .ZN(n315) );
  OR2_X1 U285 ( .A1(n616), .A2(n671), .ZN(n325) );
  AOI22_X1 U286 ( .A1(A[14]), .A2(n639), .B1(A[15]), .B2(n631), .ZN(n203) );
  OR2_X1 U287 ( .A1(n619), .A2(n667), .ZN(n326) );
  AOI22_X1 U288 ( .A1(A[23]), .A2(n640), .B1(A[24]), .B2(n578), .ZN(n223) );
  OR2_X1 U289 ( .A1(n635), .A2(n661), .ZN(n347) );
  OR2_X1 U290 ( .A1(n657), .A2(n620), .ZN(n348) );
  AOI22_X1 U291 ( .A1(A[5]), .A2(n640), .B1(A[6]), .B2(n578), .ZN(n233) );
  OR2_X1 U292 ( .A1(n619), .A2(n678), .ZN(n295) );
  AOI22_X1 U293 ( .A1(A[16]), .A2(n638), .B1(n632), .B2(A[17]), .ZN(n217) );
  OR2_X1 U294 ( .A1(n618), .A2(n665), .ZN(n359) );
  AOI22_X1 U295 ( .A1(A[20]), .A2(n638), .B1(A[21]), .B2(n613), .ZN(n216) );
  OR2_X1 U296 ( .A1(n622), .A2(n661), .ZN(n366) );
  AOI22_X1 U297 ( .A1(A[28]), .A2(n638), .B1(A[29]), .B2(n613), .ZN(n209) );
  OR2_X1 U298 ( .A1(n650), .A2(n617), .ZN(n343) );
  OR2_X1 U299 ( .A1(n623), .A2(n680), .ZN(n280) );
  AOI22_X1 U300 ( .A1(n640), .A2(A[25]), .B1(A[26]), .B2(n630), .ZN(n235) );
  AOI21_X1 U301 ( .B1(n250), .B2(n694), .A(SH[5]), .ZN(n218) );
  NAND4_X1 U302 ( .A1(n251), .A2(n252), .A3(n253), .A4(n254), .ZN(n250) );
  AOI22_X1 U303 ( .A1(A[13]), .A2(n639), .B1(A[14]), .B2(n578), .ZN(n230) );
  AOI22_X1 U304 ( .A1(A[22]), .A2(n639), .B1(A[23]), .B2(n630), .ZN(n204) );
  OAI221_X1 U305 ( .B1(n616), .B2(n659), .C1(n656), .C2(n620), .A(n573), .ZN(
        n161) );
  AOI22_X1 U306 ( .A1(A[24]), .A2(n638), .B1(A[25]), .B2(n631), .ZN(n214) );
  AOI22_X1 U307 ( .A1(A[11]), .A2(n640), .B1(A[12]), .B2(n630), .ZN(n224) );
  NAND2_X1 U308 ( .A1(SH[3]), .A2(n228), .ZN(n137) );
  NAND3_X1 U309 ( .A1(n354), .A2(n355), .A3(n226), .ZN(n173) );
  AOI22_X1 U310 ( .A1(A[15]), .A2(n640), .B1(A[16]), .B2(n630), .ZN(n226) );
  NAND3_X1 U311 ( .A1(n317), .A2(n318), .A3(n221), .ZN(n168) );
  AOI22_X1 U312 ( .A1(A[27]), .A2(n639), .B1(A[28]), .B2(n613), .ZN(n221) );
  OR2_X1 U313 ( .A1(n652), .A2(n621), .ZN(n318) );
  NAND2_X1 U314 ( .A1(SH[2]), .A2(n228), .ZN(n196) );
  NAND2_X1 U315 ( .A1(n636), .A2(A[1]), .ZN(n350) );
  OR2_X1 U316 ( .A1(n617), .A2(n682), .ZN(n351) );
  NAND3_X1 U317 ( .A1(n331), .A2(n332), .A3(n210), .ZN(n166) );
  AOI22_X1 U318 ( .A1(A[8]), .A2(n639), .B1(A[9]), .B2(n613), .ZN(n210) );
  NAND2_X1 U319 ( .A1(n344), .A2(SH[0]), .ZN(n240) );
  NOR2_X1 U320 ( .A1(n505), .A2(n506), .ZN(n245) );
  AND3_X1 U321 ( .A1(n362), .A2(n363), .A3(n364), .ZN(n125) );
  NAND2_X1 U322 ( .A1(n630), .A2(A[31]), .ZN(n362) );
  NAND2_X1 U323 ( .A1(n639), .A2(A[30]), .ZN(n363) );
  INV_X1 U324 ( .A(A[31]), .ZN(n646) );
  INV_X1 U325 ( .A(A[23]), .ZN(n659) );
  INV_X1 U326 ( .A(A[6]), .ZN(n680) );
  INV_X1 U327 ( .A(A[28]), .ZN(n653) );
  INV_X1 U328 ( .A(A[26]), .ZN(n656) );
  INV_X1 U329 ( .A(A[19]), .ZN(n664) );
  INV_X1 U330 ( .A(A[17]), .ZN(n666) );
  INV_X1 U331 ( .A(A[16]), .ZN(n667) );
  INV_X1 U332 ( .A(A[9]), .ZN(n676) );
  INV_X1 U333 ( .A(A[22]), .ZN(n661) );
  INV_X1 U334 ( .A(A[13]), .ZN(n671) );
  INV_X1 U335 ( .A(A[18]), .ZN(n665) );
  INV_X1 U336 ( .A(A[20]), .ZN(n663) );
  INV_X1 U337 ( .A(A[25]), .ZN(n657) );
  INV_X1 U338 ( .A(A[5]), .ZN(n681) );
  INV_X1 U339 ( .A(A[27]), .ZN(n654) );
  INV_X1 U340 ( .A(A[30]), .ZN(n650) );
  INV_X1 U341 ( .A(A[8]), .ZN(n677) );
  INV_X1 U342 ( .A(A[7]), .ZN(n678) );
  INV_X1 U343 ( .A(A[21]), .ZN(n662) );
  INV_X1 U344 ( .A(A[24]), .ZN(n658) );
  INV_X1 U345 ( .A(A[14]), .ZN(n670) );
  INV_X1 U346 ( .A(A[12]), .ZN(n672) );
  INV_X1 U347 ( .A(A[11]), .ZN(n673) );
  INV_X1 U348 ( .A(A[0]), .ZN(n689) );
  INV_X1 U349 ( .A(A[15]), .ZN(n669) );
  INV_X1 U350 ( .A(A[29]), .ZN(n652) );
  INV_X1 U351 ( .A(A[3]), .ZN(n684) );
  AND3_X1 U352 ( .A1(n248), .A2(SH[27]), .A3(n309), .ZN(n243) );
  OAI22_X1 U353 ( .A1(n688), .A2(n104), .B1(n107), .B2(n181), .ZN(B[1]) );
  NAND2_X1 U354 ( .A1(n154), .A2(n625), .ZN(n489) );
  NAND2_X1 U355 ( .A1(n154), .A2(n642), .ZN(n482) );
  INV_X1 U356 ( .A(A[2]), .ZN(n685) );
  AOI22_X1 U357 ( .A1(A[2]), .A2(n638), .B1(A[3]), .B2(n613), .ZN(n197) );
  AOI22_X1 U358 ( .A1(A[4]), .A2(n639), .B1(A[5]), .B2(n632), .ZN(n212) );
  AOI22_X1 U359 ( .A1(A[3]), .A2(n640), .B1(A[4]), .B2(n632), .ZN(n220) );
  INV_X1 U360 ( .A(A[4]), .ZN(n682) );
  AOI22_X1 U361 ( .A1(A[10]), .A2(n640), .B1(A[11]), .B2(n631), .ZN(n199) );
  AOI22_X1 U362 ( .A1(A[9]), .A2(n640), .B1(A[10]), .B2(n632), .ZN(n232) );
  INV_X1 U363 ( .A(A[10]), .ZN(n675) );
  OAI221_X1 U364 ( .B1(n594), .B2(n689), .C1(n620), .C2(n684), .A(n231), .ZN(
        n153) );
  AOI22_X1 U365 ( .A1(A[1]), .A2(n639), .B1(A[2]), .B2(n631), .ZN(n231) );
  NAND2_X1 U366 ( .A1(n604), .A2(n584), .ZN(n616) );
  INV_X1 U367 ( .A(n637), .ZN(n635) );
  OAI221_X1 U368 ( .B1(n133), .B2(n692), .C1(n134), .C2(n693), .A(n135), .ZN(
        B[27]) );
  OAI22_X1 U369 ( .A1(n189), .A2(n690), .B1(n190), .B2(n693), .ZN(B[16]) );
  OAI22_X1 U370 ( .A1(n645), .A2(n112), .B1(n113), .B2(n114), .ZN(B[31]) );
  INV_X1 U371 ( .A(n624), .ZN(n617) );
  INV_X1 U372 ( .A(n599), .ZN(n618) );
  INV_X1 U374 ( .A(n624), .ZN(n619) );
  INV_X1 U375 ( .A(n597), .ZN(n620) );
  INV_X1 U376 ( .A(n597), .ZN(n621) );
  INV_X1 U377 ( .A(n599), .ZN(n622) );
  INV_X1 U378 ( .A(n598), .ZN(n623) );
  NOR3_X1 U379 ( .A1(n329), .A2(n330), .A3(n660), .ZN(n92) );
  INV_X1 U380 ( .A(n572), .ZN(n683) );
  AOI22_X1 U381 ( .A1(n587), .A2(n628), .B1(n572), .B2(n642), .ZN(n91) );
  NAND2_X1 U382 ( .A1(n636), .A2(A[29]), .ZN(n364) );
  NAND4_X1 U383 ( .A1(n244), .A2(n243), .A3(n245), .A4(n610), .ZN(n283) );
  NAND4_X1 U384 ( .A1(n242), .A2(n244), .A3(n245), .A4(n243), .ZN(n241) );
  AND3_X1 U385 ( .A1(SH[18]), .A2(SH[17]), .A3(SH[19]), .ZN(n247) );
  NAND2_X1 U386 ( .A1(n241), .A2(SH[31]), .ZN(n344) );
  NAND2_X1 U387 ( .A1(SH[31]), .A2(n283), .ZN(n228) );
  INV_X1 U388 ( .A(SH[31]), .ZN(n694) );
  AND2_X1 U389 ( .A1(n136), .A2(n696), .ZN(n376) );
  NOR2_X1 U390 ( .A1(n196), .A2(n696), .ZN(n387) );
  NOR2_X1 U391 ( .A1(n697), .A2(n137), .ZN(n261) );
  INV_X1 U392 ( .A(n137), .ZN(n696) );
  AOI222_X1 U393 ( .A1(n600), .A2(n643), .B1(n686), .B2(n626), .C1(n586), .C2(
        n628), .ZN(n133) );
  AOI22_X1 U394 ( .A1(n600), .A2(n633), .B1(n629), .B2(n592), .ZN(n184) );
  AOI22_X1 U395 ( .A1(n598), .A2(A[1]), .B1(n632), .B2(A[0]), .ZN(n121) );
  NOR2_X1 U396 ( .A1(n604), .A2(n383), .ZN(n272) );
  INV_X1 U397 ( .A(n383), .ZN(n698) );
  AOI22_X1 U398 ( .A1(n633), .A2(n603), .B1(n629), .B2(n145), .ZN(n188) );
  AOI222_X1 U399 ( .A1(n603), .A2(n643), .B1(n627), .B2(n143), .C1(n144), .C2(
        n628), .ZN(n88) );
  OAI222_X1 U400 ( .A1(n388), .A2(n690), .B1(n645), .B2(n191), .C1(n352), .C2(
        n693), .ZN(B[15]) );
  OR2_X1 U401 ( .A1(n616), .A2(n662), .ZN(n290) );
  OR2_X1 U402 ( .A1(n635), .A2(n682), .ZN(n294) );
  OR2_X1 U403 ( .A1(n596), .A2(n676), .ZN(n305) );
  OR2_X1 U404 ( .A1(n616), .A2(n677), .ZN(n314) );
  OR2_X1 U405 ( .A1(n596), .A2(n658), .ZN(n367) );
  OR2_X1 U406 ( .A1(n594), .A2(n657), .ZN(n371) );
  OR2_X1 U407 ( .A1(n616), .A2(n663), .ZN(n302) );
  OR2_X1 U408 ( .A1(n616), .A2(n681), .ZN(n286) );
  OR2_X1 U409 ( .A1(n596), .A2(n684), .ZN(n279) );
  OR2_X1 U410 ( .A1(n594), .A2(n656), .ZN(n317) );
  OR2_X1 U411 ( .A1(n594), .A2(n673), .ZN(n379) );
  OR2_X1 U412 ( .A1(n596), .A2(n664), .ZN(n365) );
  OR2_X1 U413 ( .A1(n616), .A2(n672), .ZN(n335) );
  OR2_X1 U414 ( .A1(n596), .A2(n654), .ZN(n342) );
  OR2_X1 U415 ( .A1(n594), .A2(n669), .ZN(n358) );
  AOI22_X1 U416 ( .A1(n634), .A2(n173), .B1(n629), .B2(n168), .ZN(n195) );
  OAI22_X1 U417 ( .A1(n117), .A2(n112), .B1(n113), .B2(n118), .ZN(B[30]) );
  OR2_X1 U418 ( .A1(n618), .A2(n666), .ZN(n355) );
  OR2_X1 U419 ( .A1(n616), .A2(n670), .ZN(n354) );
  OAI222_X1 U420 ( .A1(n127), .A2(n690), .B1(n125), .B2(n191), .C1(n322), .C2(
        n693), .ZN(B[13]) );
  AOI222_X1 U421 ( .A1(n148), .A2(n629), .B1(n144), .B2(n642), .C1(n137), .C2(
        n101), .ZN(n322) );
  OR3_X1 U422 ( .A1(SH[14]), .A2(SH[15]), .A3(SH[13]), .ZN(n258) );
  OR2_X1 U423 ( .A1(n596), .A2(n678), .ZN(n331) );
  OR2_X1 U424 ( .A1(n621), .A2(n675), .ZN(n332) );
  NOR4_X1 U425 ( .A1(n257), .A2(SH[16]), .A3(SH[18]), .A4(n593), .ZN(n252) );
  OR3_X1 U426 ( .A1(SH[20]), .A2(SH[21]), .A3(SH[19]), .ZN(n257) );
  OR3_X1 U427 ( .A1(SH[26]), .A2(SH[27]), .A3(SH[25]), .ZN(n256) );
  OAI221_X1 U428 ( .B1(n134), .B2(n690), .C1(n133), .C2(n693), .A(n208), .ZN(
        B[11]) );
  INV_X1 U429 ( .A(n213), .ZN(n655) );
  AND3_X1 U430 ( .A1(SH[24]), .A2(SH[23]), .A3(SH[25]), .ZN(n248) );
  NOR4_X1 U431 ( .A1(n258), .A2(SH[10]), .A3(SH[12]), .A4(SH[11]), .ZN(n251)
         );
  NAND4_X1 U432 ( .A1(SH[10]), .A2(SH[12]), .A3(SH[11]), .A4(SH[13]), .ZN(n505) );
  OR4_X1 U433 ( .A1(SH[6]), .A2(SH[7]), .A3(SH[8]), .A4(SH[9]), .ZN(n255) );
  AND3_X1 U434 ( .A1(SH[30]), .A2(SH[29]), .A3(SH[6]), .ZN(n249) );
  NOR4_X1 U435 ( .A1(n255), .A2(n611), .A3(SH[30]), .A4(SH[29]), .ZN(n254) );
  AND2_X1 U436 ( .A1(SH[28]), .A2(SH[26]), .ZN(n309) );
  AOI221_X1 U437 ( .B1(n167), .B2(n626), .C1(n583), .C2(n641), .A(n649), .ZN(
        n388) );
  AND2_X1 U438 ( .A1(n167), .A2(n627), .ZN(n356) );
  AND2_X1 U439 ( .A1(n167), .A2(n634), .ZN(n374) );
  AOI22_X1 U440 ( .A1(n634), .A2(n586), .B1(n629), .B2(n167), .ZN(n165) );
  NOR4_X1 U441 ( .A1(n256), .A2(SH[22]), .A3(SH[24]), .A4(SH[23]), .ZN(n253)
         );
  INV_X1 U442 ( .A(n615), .ZN(n629) );
  INV_X1 U443 ( .A(n595), .ZN(n636) );
  INV_X1 U444 ( .A(n595), .ZN(n637) );
endmodule


module SHIFTER_M32_N5 ( A, B, LEFT_RIGHT, OUTPUT );
  input [31:0] A;
  input [31:0] B;
  output [31:0] OUTPUT;
  input LEFT_RIGHT;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, n42, n44, n49, n50, n52, n53, n57,
         n58, n59, n61, n63, n64, n67, n68, n70, n71, n72, n73, net131953,
         net131968, net131973, net131978, net133051, net133049, net133047,
         net133045, net133043, net133041, net133037, net133033, net133065,
         n140, n142, n143, n144, n145, n146, n147;
  assign OUTPUT[5] = net131953;
  assign OUTPUT[3] = net131968;
  assign OUTPUT[31] = net131973;
  assign OUTPUT[4] = net131978;

  SHIFTER_M32_N5_DW01_ash_0 sll_29 ( .A(A), .DATA_TC(1'b0), .SH(B), .SH_TC(
        1'b1), .B({N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, 
        N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37, N36, N35, N34}) );
  SHIFTER_M32_N5_DW_rash_0 srl_27 ( .A(A), .DATA_TC(1'b0), .SH(B), .SH_TC(1'b1), .B({N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
        N4, N3, N2}) );
  MUX2_X1 U1 ( .A(N47), .B(N15), .S(net133033), .Z(OUTPUT[13]) );
  INV_X1 U2 ( .A(N10), .ZN(n140) );
  NAND2_X1 U7 ( .A1(n142), .A2(n143), .ZN(OUTPUT[8]) );
  OR2_X1 U8 ( .A1(n144), .A2(n140), .ZN(n142) );
  NAND2_X1 U9 ( .A1(net133043), .A2(N42), .ZN(n143) );
  MUX2_X1 U10 ( .A(N55), .B(N23), .S(net133033), .Z(OUTPUT[21]) );
  MUX2_X1 U11 ( .A(N38), .B(N6), .S(net133033), .Z(net131978) );
  MUX2_X1 U12 ( .A(N5), .B(N37), .S(LEFT_RIGHT), .Z(net131968) );
  MUX2_X1 U13 ( .A(N27), .B(N59), .S(LEFT_RIGHT), .Z(OUTPUT[25]) );
  MUX2_X1 U14 ( .A(N29), .B(N61), .S(LEFT_RIGHT), .Z(OUTPUT[27]) );
  MUX2_X1 U15 ( .A(N7), .B(N39), .S(LEFT_RIGHT), .Z(net131953) );
  MUX2_X1 U16 ( .A(N8), .B(N40), .S(LEFT_RIGHT), .Z(OUTPUT[6]) );
  MUX2_X1 U17 ( .A(N28), .B(N60), .S(LEFT_RIGHT), .Z(OUTPUT[26]) );
  MUX2_X1 U18 ( .A(N18), .B(N50), .S(LEFT_RIGHT), .Z(OUTPUT[16]) );
  MUX2_X1 U19 ( .A(N19), .B(N51), .S(LEFT_RIGHT), .Z(OUTPUT[17]) );
  MUX2_X1 U20 ( .A(N4), .B(N36), .S(LEFT_RIGHT), .Z(OUTPUT[2]) );
  MUX2_X1 U21 ( .A(N3), .B(N35), .S(LEFT_RIGHT), .Z(OUTPUT[1]) );
  BUF_X1 U22 ( .A(n146), .Z(n144) );
  AOI22_X1 U23 ( .A1(N33), .A2(net133033), .B1(N65), .B2(n144), .ZN(n49) );
  BUF_X1 U24 ( .A(LEFT_RIGHT), .Z(n146) );
  BUF_X1 U25 ( .A(n146), .Z(net133041) );
  BUF_X1 U26 ( .A(n146), .Z(net133037) );
  BUF_X1 U27 ( .A(n147), .Z(n145) );
  INV_X1 U28 ( .A(n145), .ZN(net133033) );
  BUF_X1 U29 ( .A(LEFT_RIGHT), .Z(n147) );
  BUF_X1 U30 ( .A(n147), .Z(net133049) );
  BUF_X1 U31 ( .A(n147), .Z(net133051) );
  BUF_X1 U32 ( .A(LEFT_RIGHT), .Z(net133065) );
  BUF_X1 U33 ( .A(net133065), .Z(net133045) );
  BUF_X1 U34 ( .A(net133065), .Z(net133047) );
  BUF_X1 U35 ( .A(net133065), .Z(net133043) );
  AOI22_X1 U36 ( .A1(N25), .A2(net133033), .B1(N57), .B2(net133045), .ZN(n58)
         );
  INV_X1 U37 ( .A(n44), .ZN(OUTPUT[7]) );
  INV_X1 U38 ( .A(n49), .ZN(net131973) );
  INV_X1 U39 ( .A(n58), .ZN(OUTPUT[23]) );
  INV_X1 U40 ( .A(n68), .ZN(OUTPUT[14]) );
  INV_X1 U41 ( .A(n63), .ZN(OUTPUT[19]) );
  AOI22_X1 U42 ( .A1(N24), .A2(net133033), .B1(N56), .B2(net133045), .ZN(n59)
         );
  AOI22_X1 U43 ( .A1(N30), .A2(net133033), .B1(N62), .B2(net133041), .ZN(n53)
         );
  AOI22_X1 U44 ( .A1(N16), .A2(net133033), .B1(N48), .B2(net133049), .ZN(n68)
         );
  AOI22_X1 U45 ( .A1(N22), .A2(net133033), .B1(N54), .B2(net133045), .ZN(n61)
         );
  AOI22_X1 U46 ( .A1(N20), .A2(net133033), .B1(N52), .B2(net133047), .ZN(n64)
         );
  AOI22_X1 U47 ( .A1(N21), .A2(net133033), .B1(N53), .B2(net133047), .ZN(n63)
         );
  INV_X1 U48 ( .A(n61), .ZN(OUTPUT[20]) );
  AOI22_X1 U49 ( .A1(N13), .A2(net133033), .B1(N45), .B2(net133051), .ZN(n71)
         );
  INV_X1 U50 ( .A(n52), .ZN(OUTPUT[29]) );
  AOI22_X1 U51 ( .A1(N14), .A2(net133033), .B1(N46), .B2(net133051), .ZN(n70)
         );
  AOI22_X1 U52 ( .A1(N17), .A2(net133033), .B1(N49), .B2(net133049), .ZN(n67)
         );
  INV_X1 U53 ( .A(n67), .ZN(OUTPUT[15]) );
  INV_X1 U54 ( .A(n42), .ZN(OUTPUT[9]) );
  AOI22_X1 U55 ( .A1(N11), .A2(net133033), .B1(N43), .B2(net133037), .ZN(n42)
         );
  INV_X1 U56 ( .A(n59), .ZN(OUTPUT[22]) );
  AOI22_X1 U57 ( .A1(N32), .A2(net133033), .B1(N64), .B2(net133041), .ZN(n50)
         );
  INV_X1 U58 ( .A(n72), .ZN(OUTPUT[10]) );
  INV_X1 U59 ( .A(n57), .ZN(OUTPUT[24]) );
  INV_X1 U60 ( .A(n71), .ZN(OUTPUT[11]) );
  INV_X1 U61 ( .A(n64), .ZN(OUTPUT[18]) );
  INV_X1 U62 ( .A(n50), .ZN(OUTPUT[30]) );
  AOI22_X1 U63 ( .A1(N26), .A2(net133033), .B1(N58), .B2(net133043), .ZN(n57)
         );
  AOI22_X1 U64 ( .A1(N12), .A2(net133033), .B1(N44), .B2(net133051), .ZN(n72)
         );
  INV_X1 U65 ( .A(n70), .ZN(OUTPUT[12]) );
  AOI22_X1 U66 ( .A1(N2), .A2(net133033), .B1(N34), .B2(net133051), .ZN(n73)
         );
  AOI22_X1 U67 ( .A1(N9), .A2(net133033), .B1(N41), .B2(net133037), .ZN(n44)
         );
  INV_X1 U68 ( .A(n73), .ZN(OUTPUT[0]) );
  INV_X1 U69 ( .A(n53), .ZN(OUTPUT[28]) );
  AOI22_X1 U70 ( .A1(N31), .A2(net133033), .B1(N63), .B2(net133041), .ZN(n52)
         );
endmodule


module PGnet_0 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_30 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_29 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_28 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_27 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_26 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_25 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_24 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_23 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_22 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_21 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_20 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_19 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_18 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_17 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_16 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_15 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_14 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_13 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_12 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_11 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_10 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_9 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_8 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_7 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_6 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_5 ( A, B, p, g );
  input A, B;
  output p, g;
  wire   n1;

  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  CLKBUF_X1 U1 ( .A(B), .Z(n1) );
  AND2_X1 U3 ( .A1(n1), .A2(A), .ZN(g) );
endmodule


module PGnet_4 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_3 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_2 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PGnet_1 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module G_0 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n2) );
endmodule


module G_9 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
endmodule


module PG_0 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n2;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n2), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(p1), .B2(g2), .A(g1), .ZN(n2) );
endmodule


module PG_26 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_25 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_24 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_23 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n7), .B2(n8), .A(n9), .ZN(g_Out) );
  INV_X1 U2 ( .A(g2), .ZN(n7) );
  INV_X1 U3 ( .A(p1), .ZN(n8) );
  INV_X1 U4 ( .A(g1), .ZN(n9) );
  AND2_X1 U5 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_22 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
endmodule


module PG_21 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n7), .B2(n8), .A(n9), .ZN(g_Out) );
  INV_X1 U2 ( .A(g2), .ZN(n7) );
  INV_X1 U3 ( .A(p1), .ZN(n8) );
  INV_X1 U4 ( .A(g1), .ZN(n9) );
  AND2_X1 U5 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_20 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_19 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_18 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_17 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
endmodule


module PG_16 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_15 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_14 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
endmodule


module PG_13 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
endmodule


module G_8 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
endmodule


module PG_12 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
endmodule


module PG_11 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_10 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_9 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_8 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_7 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_6 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module G_7 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
endmodule


module PG_5 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(p_Out) );
endmodule


module PG_4 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  AOI21_X1 U1 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U3 ( .A(n8), .ZN(g_Out) );
endmodule


module PG_3 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U2 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
endmodule


module G_6 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
endmodule


module G_5 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X2 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
endmodule


module PG_2 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  AOI21_X1 U1 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  INV_X1 U3 ( .A(n8), .ZN(g_Out) );
endmodule


module PG_1 ( p1, g1, p2, g2, p_Out, g_Out );
  input p1, g1, p2, g2;
  output p_Out, g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(p_Out) );
  AOI21_X1 U3 ( .B1(g2), .B2(p1), .A(g1), .ZN(n8) );
endmodule


module G_4 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
endmodule


module G_3 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
endmodule


module G_2 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
endmodule


module G_1 ( p1, g1, g2, g_Out );
  input p1, g1, g2;
  output g_Out;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(g_Out) );
  AOI21_X1 U2 ( .B1(p1), .B2(g2), .A(g1), .ZN(n8) );
endmodule


module Cg ( A, B, cin0, cout );
  input [31:0] A;
  input [31:0] B;
  output [7:0] cout;
  input cin0;
  wire   n3, n6, n7, p0, g0, \gsignal[4][31] , \gsignal[4][27] ,
         \gsignal[3][31] , \gsignal[3][23] , \gsignal[3][15] ,
         \gsignal[2][31] , \gsignal[2][27] , \gsignal[2][23] ,
         \gsignal[2][19] , \gsignal[2][15] , \gsignal[2][11] , \gsignal[2][7] ,
         \gsignal[1][31] , \gsignal[1][29] , \gsignal[1][27] ,
         \gsignal[1][25] , \gsignal[1][23] , \gsignal[1][21] ,
         \gsignal[1][19] , \gsignal[1][17] , \gsignal[1][15] ,
         \gsignal[1][13] , \gsignal[1][11] , \gsignal[1][9] , \gsignal[1][7] ,
         \gsignal[1][5] , \gsignal[1][3] , \gsignal[1][1] , \gsignal[0][31] ,
         \gsignal[0][30] , \gsignal[0][29] , \gsignal[0][28] ,
         \gsignal[0][27] , \gsignal[0][26] , \gsignal[0][25] ,
         \gsignal[0][24] , \gsignal[0][23] , \gsignal[0][22] ,
         \gsignal[0][21] , \gsignal[0][20] , \gsignal[0][19] ,
         \gsignal[0][18] , \gsignal[0][17] , \gsignal[0][16] ,
         \gsignal[0][15] , \gsignal[0][14] , \gsignal[0][13] ,
         \gsignal[0][12] , \gsignal[0][11] , \gsignal[0][10] , \gsignal[0][9] ,
         \gsignal[0][8] , \gsignal[0][7] , \gsignal[0][6] , \gsignal[0][5] ,
         \gsignal[0][4] , \gsignal[0][3] , \gsignal[0][2] , \gsignal[0][1] ,
         \gsignal[0][0] , \psignal[4][31] , \psignal[4][27] , \psignal[3][31] ,
         \psignal[3][23] , \psignal[3][15] , \psignal[2][31] ,
         \psignal[2][27] , \psignal[2][23] , \psignal[2][19] ,
         \psignal[2][15] , \psignal[2][11] , \psignal[2][7] , \psignal[1][31] ,
         \psignal[1][29] , \psignal[1][27] , \psignal[1][25] ,
         \psignal[1][23] , \psignal[1][21] , \psignal[1][19] ,
         \psignal[1][17] , \psignal[1][15] , \psignal[1][13] ,
         \psignal[1][11] , \psignal[1][9] , \psignal[1][7] , \psignal[1][5] ,
         \psignal[1][3] , \psignal[0][31] , \psignal[0][30] , \psignal[0][29] ,
         \psignal[0][28] , \psignal[0][27] , \psignal[0][26] ,
         \psignal[0][25] , \psignal[0][24] , \psignal[0][23] ,
         \psignal[0][22] , \psignal[0][21] , \psignal[0][20] ,
         \psignal[0][19] , \psignal[0][18] , \psignal[0][17] ,
         \psignal[0][16] , \psignal[0][15] , \psignal[0][14] ,
         \psignal[0][13] , \psignal[0][12] , \psignal[0][11] ,
         \psignal[0][10] , \psignal[0][9] , \psignal[0][8] , \psignal[0][7] ,
         \psignal[0][6] , \psignal[0][5] , \psignal[0][4] , \psignal[0][3] ,
         \psignal[0][2] , \psignal[0][1] ;
  assign cout[3] = n3;

  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(p0) );
  PGnet_0 PGN1_31 ( .A(A[31]), .B(B[31]), .p(\psignal[0][31] ), .g(
        \gsignal[0][31] ) );
  PGnet_30 PGN1_30 ( .A(A[30]), .B(B[30]), .p(\psignal[0][30] ), .g(
        \gsignal[0][30] ) );
  PGnet_29 PGN1_29 ( .A(A[29]), .B(B[29]), .p(\psignal[0][29] ), .g(
        \gsignal[0][29] ) );
  PGnet_28 PGN1_28 ( .A(A[28]), .B(B[28]), .p(\psignal[0][28] ), .g(
        \gsignal[0][28] ) );
  PGnet_27 PGN1_27 ( .A(A[27]), .B(B[27]), .p(\psignal[0][27] ), .g(
        \gsignal[0][27] ) );
  PGnet_26 PGN1_26 ( .A(A[26]), .B(B[26]), .p(\psignal[0][26] ), .g(
        \gsignal[0][26] ) );
  PGnet_25 PGN1_25 ( .A(A[25]), .B(B[25]), .p(\psignal[0][25] ), .g(
        \gsignal[0][25] ) );
  PGnet_24 PGN1_24 ( .A(A[24]), .B(B[24]), .p(\psignal[0][24] ), .g(
        \gsignal[0][24] ) );
  PGnet_23 PGN1_23 ( .A(A[23]), .B(B[23]), .p(\psignal[0][23] ), .g(
        \gsignal[0][23] ) );
  PGnet_22 PGN1_22 ( .A(A[22]), .B(B[22]), .p(\psignal[0][22] ), .g(
        \gsignal[0][22] ) );
  PGnet_21 PGN1_21 ( .A(A[21]), .B(B[21]), .p(\psignal[0][21] ), .g(
        \gsignal[0][21] ) );
  PGnet_20 PGN1_20 ( .A(A[20]), .B(B[20]), .p(\psignal[0][20] ), .g(
        \gsignal[0][20] ) );
  PGnet_19 PGN1_19 ( .A(A[19]), .B(B[19]), .p(\psignal[0][19] ), .g(
        \gsignal[0][19] ) );
  PGnet_18 PGN1_18 ( .A(A[18]), .B(B[18]), .p(\psignal[0][18] ), .g(
        \gsignal[0][18] ) );
  PGnet_17 PGN1_17 ( .A(A[17]), .B(B[17]), .p(\psignal[0][17] ), .g(
        \gsignal[0][17] ) );
  PGnet_16 PGN1_16 ( .A(A[16]), .B(B[16]), .p(\psignal[0][16] ), .g(
        \gsignal[0][16] ) );
  PGnet_15 PGN1_15 ( .A(A[15]), .B(B[15]), .p(\psignal[0][15] ), .g(
        \gsignal[0][15] ) );
  PGnet_14 PGN1_14 ( .A(A[14]), .B(B[14]), .p(\psignal[0][14] ), .g(
        \gsignal[0][14] ) );
  PGnet_13 PGN1_13 ( .A(A[13]), .B(B[13]), .p(\psignal[0][13] ), .g(
        \gsignal[0][13] ) );
  PGnet_12 PGN1_12 ( .A(A[12]), .B(B[12]), .p(\psignal[0][12] ), .g(
        \gsignal[0][12] ) );
  PGnet_11 PGN1_11 ( .A(A[11]), .B(B[11]), .p(\psignal[0][11] ), .g(
        \gsignal[0][11] ) );
  PGnet_10 PGN1_10 ( .A(A[10]), .B(B[10]), .p(\psignal[0][10] ), .g(
        \gsignal[0][10] ) );
  PGnet_9 PGN1_9 ( .A(A[9]), .B(B[9]), .p(\psignal[0][9] ), .g(\gsignal[0][9] ) );
  PGnet_8 PGN1_8 ( .A(A[8]), .B(B[8]), .p(\psignal[0][8] ), .g(\gsignal[0][8] ) );
  PGnet_7 PGN1_7 ( .A(A[7]), .B(B[7]), .p(\psignal[0][7] ), .g(\gsignal[0][7] ) );
  PGnet_6 PGN1_6 ( .A(A[6]), .B(B[6]), .p(\psignal[0][6] ), .g(\gsignal[0][6] ) );
  PGnet_5 PGN1_5 ( .A(A[5]), .B(B[5]), .p(\psignal[0][5] ), .g(\gsignal[0][5] ) );
  PGnet_4 PGN1_4 ( .A(A[4]), .B(B[4]), .p(\psignal[0][4] ), .g(\gsignal[0][4] ) );
  PGnet_3 PGN1_3 ( .A(A[3]), .B(B[3]), .p(\psignal[0][3] ), .g(\gsignal[0][3] ) );
  PGnet_2 PGN1_2 ( .A(A[2]), .B(B[2]), .p(\psignal[0][2] ), .g(\gsignal[0][2] ) );
  PGnet_1 PGN1_1 ( .A(A[1]), .B(B[1]), .p(\psignal[0][1] ), .g(\gsignal[0][1] ) );
  G_0 PGN0_0 ( .p1(p0), .g1(g0), .g2(cin0), .g_Out(\gsignal[0][0] ) );
  G_9 g0_0_1 ( .p1(\psignal[0][1] ), .g1(\gsignal[0][1] ), .g2(\gsignal[0][0] ), .g_Out(\gsignal[1][1] ) );
  PG_0 PGelements_0_3 ( .p1(\psignal[0][3] ), .g1(\gsignal[0][3] ), .p2(
        \psignal[0][2] ), .g2(\gsignal[0][2] ), .p_Out(\psignal[1][3] ), 
        .g_Out(\gsignal[1][3] ) );
  PG_26 PGelements_0_5 ( .p1(\psignal[0][5] ), .g1(\gsignal[0][5] ), .p2(
        \psignal[0][4] ), .g2(\gsignal[0][4] ), .p_Out(\psignal[1][5] ), 
        .g_Out(\gsignal[1][5] ) );
  PG_25 PGelements_0_7 ( .p1(\psignal[0][7] ), .g1(\gsignal[0][7] ), .p2(
        \psignal[0][6] ), .g2(\gsignal[0][6] ), .p_Out(\psignal[1][7] ), 
        .g_Out(\gsignal[1][7] ) );
  PG_24 PGelements_0_9 ( .p1(\psignal[0][9] ), .g1(\gsignal[0][9] ), .p2(
        \psignal[0][8] ), .g2(\gsignal[0][8] ), .p_Out(\psignal[1][9] ), 
        .g_Out(\gsignal[1][9] ) );
  PG_23 PGelements_0_11 ( .p1(\psignal[0][11] ), .g1(\gsignal[0][11] ), .p2(
        \psignal[0][10] ), .g2(\gsignal[0][10] ), .p_Out(\psignal[1][11] ), 
        .g_Out(\gsignal[1][11] ) );
  PG_22 PGelements_0_13 ( .p1(\psignal[0][13] ), .g1(\gsignal[0][13] ), .p2(
        \psignal[0][12] ), .g2(\gsignal[0][12] ), .p_Out(\psignal[1][13] ), 
        .g_Out(\gsignal[1][13] ) );
  PG_21 PGelements_0_15 ( .p1(\psignal[0][15] ), .g1(\gsignal[0][15] ), .p2(
        \psignal[0][14] ), .g2(\gsignal[0][14] ), .p_Out(\psignal[1][15] ), 
        .g_Out(\gsignal[1][15] ) );
  PG_20 PGelements_0_17 ( .p1(\psignal[0][17] ), .g1(\gsignal[0][17] ), .p2(
        \psignal[0][16] ), .g2(\gsignal[0][16] ), .p_Out(\psignal[1][17] ), 
        .g_Out(\gsignal[1][17] ) );
  PG_19 PGelements_0_19 ( .p1(\psignal[0][19] ), .g1(\gsignal[0][19] ), .p2(
        \psignal[0][18] ), .g2(\gsignal[0][18] ), .p_Out(\psignal[1][19] ), 
        .g_Out(\gsignal[1][19] ) );
  PG_18 PGelements_0_21 ( .p1(\psignal[0][21] ), .g1(\gsignal[0][21] ), .p2(
        \psignal[0][20] ), .g2(\gsignal[0][20] ), .p_Out(\psignal[1][21] ), 
        .g_Out(\gsignal[1][21] ) );
  PG_17 PGelements_0_23 ( .p1(\psignal[0][23] ), .g1(\gsignal[0][23] ), .p2(
        \psignal[0][22] ), .g2(\gsignal[0][22] ), .p_Out(\psignal[1][23] ), 
        .g_Out(\gsignal[1][23] ) );
  PG_16 PGelements_0_25 ( .p1(\psignal[0][25] ), .g1(\gsignal[0][25] ), .p2(
        \psignal[0][24] ), .g2(\gsignal[0][24] ), .p_Out(\psignal[1][25] ), 
        .g_Out(\gsignal[1][25] ) );
  PG_15 PGelements_0_27 ( .p1(\psignal[0][27] ), .g1(\gsignal[0][27] ), .p2(
        \psignal[0][26] ), .g2(\gsignal[0][26] ), .p_Out(\psignal[1][27] ), 
        .g_Out(\gsignal[1][27] ) );
  PG_14 PGelements_0_29 ( .p1(\psignal[0][29] ), .g1(\gsignal[0][29] ), .p2(
        \psignal[0][28] ), .g2(\gsignal[0][28] ), .p_Out(\psignal[1][29] ), 
        .g_Out(\gsignal[1][29] ) );
  PG_13 PGelements_0_31 ( .p1(\psignal[0][31] ), .g1(\gsignal[0][31] ), .p2(
        \psignal[0][30] ), .g2(\gsignal[0][30] ), .p_Out(\psignal[1][31] ), 
        .g_Out(\gsignal[1][31] ) );
  G_8 g0_1_3 ( .p1(\psignal[1][3] ), .g1(\gsignal[1][3] ), .g2(\gsignal[1][1] ), .g_Out(n7) );
  PG_12 PGelements_1_7 ( .p1(\psignal[1][7] ), .g1(\gsignal[1][7] ), .p2(
        \psignal[1][5] ), .g2(\gsignal[1][5] ), .p_Out(\psignal[2][7] ), 
        .g_Out(\gsignal[2][7] ) );
  PG_11 PGelements_1_11 ( .p1(\psignal[1][11] ), .g1(\gsignal[1][11] ), .p2(
        \psignal[1][9] ), .g2(\gsignal[1][9] ), .p_Out(\psignal[2][11] ), 
        .g_Out(\gsignal[2][11] ) );
  PG_10 PGelements_1_15 ( .p1(\psignal[1][15] ), .g1(\gsignal[1][15] ), .p2(
        \psignal[1][13] ), .g2(\gsignal[1][13] ), .p_Out(\psignal[2][15] ), 
        .g_Out(\gsignal[2][15] ) );
  PG_9 PGelements_1_19 ( .p1(\psignal[1][19] ), .g1(\gsignal[1][19] ), .p2(
        \psignal[1][17] ), .g2(\gsignal[1][17] ), .p_Out(\psignal[2][19] ), 
        .g_Out(\gsignal[2][19] ) );
  PG_8 PGelements_1_23 ( .p1(\psignal[1][23] ), .g1(\gsignal[1][23] ), .p2(
        \psignal[1][21] ), .g2(\gsignal[1][21] ), .p_Out(\psignal[2][23] ), 
        .g_Out(\gsignal[2][23] ) );
  PG_7 PGelements_1_27 ( .p1(\psignal[1][27] ), .g1(\gsignal[1][27] ), .p2(
        \psignal[1][25] ), .g2(\gsignal[1][25] ), .p_Out(\psignal[2][27] ), 
        .g_Out(\gsignal[2][27] ) );
  PG_6 PGelements_1_31 ( .p1(\psignal[1][31] ), .g1(\gsignal[1][31] ), .p2(
        \psignal[1][29] ), .g2(\gsignal[1][29] ), .p_Out(\psignal[2][31] ), 
        .g_Out(\gsignal[2][31] ) );
  G_7 g0_2_7 ( .p1(\psignal[2][7] ), .g1(\gsignal[2][7] ), .g2(n7), .g_Out(n6)
         );
  PG_5 PGelements_2_15 ( .p1(\psignal[2][15] ), .g1(\gsignal[2][15] ), .p2(
        \psignal[2][11] ), .g2(\gsignal[2][11] ), .p_Out(\psignal[3][15] ), 
        .g_Out(\gsignal[3][15] ) );
  PG_4 PGelements_2_23 ( .p1(\psignal[2][23] ), .g1(\gsignal[2][23] ), .p2(
        \psignal[2][19] ), .g2(\gsignal[2][19] ), .p_Out(\psignal[3][23] ), 
        .g_Out(\gsignal[3][23] ) );
  PG_3 PGelements_2_31 ( .p1(\psignal[2][31] ), .g1(\gsignal[2][31] ), .p2(
        \psignal[2][27] ), .g2(\gsignal[2][27] ), .p_Out(\psignal[3][31] ), 
        .g_Out(\gsignal[3][31] ) );
  G_6 g1_3_11 ( .p1(\psignal[2][11] ), .g1(\gsignal[2][11] ), .g2(cout[1]), 
        .g_Out(cout[2]) );
  G_5 g1_3_15 ( .p1(\psignal[3][15] ), .g1(\gsignal[3][15] ), .g2(n6), .g_Out(
        n3) );
  PG_2 pg1_3_27 ( .p1(\psignal[2][27] ), .g1(\gsignal[2][27] ), .p2(
        \psignal[3][15] ), .g2(\gsignal[3][15] ), .p_Out(\psignal[4][27] ), 
        .g_Out(\gsignal[4][27] ) );
  PG_1 pg1_3_31 ( .p1(\psignal[3][31] ), .g1(\gsignal[3][31] ), .p2(
        \psignal[3][15] ), .g2(\gsignal[3][15] ), .p_Out(\psignal[4][31] ), 
        .g_Out(\gsignal[4][31] ) );
  G_4 g1_4_19 ( .p1(\psignal[2][19] ), .g1(\gsignal[2][19] ), .g2(n3), .g_Out(
        cout[4]) );
  G_3 g1_4_23 ( .p1(\psignal[3][23] ), .g1(\gsignal[3][23] ), .g2(n3), .g_Out(
        cout[5]) );
  G_2 g1_4_27 ( .p1(\psignal[4][27] ), .g1(\gsignal[4][27] ), .g2(n3), .g_Out(
        cout[6]) );
  G_1 g1_4_31 ( .p1(\psignal[4][31] ), .g1(\gsignal[4][31] ), .g2(n3), .g_Out(
        cout[7]) );
  BUF_X1 U1 ( .A(n7), .Z(cout[0]) );
  BUF_X2 U3 ( .A(n6), .Z(cout[1]) );
  AND2_X1 U4 ( .A1(B[0]), .A2(A[0]), .ZN(g0) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U1 ( .A(n2), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n3), .B2(Ci), .ZN(n2) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_0 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n6, n7, n8, n9, n18;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(n6), .ZN(s[3]) );
  AOI22_X1 U4 ( .A1(out0[3]), .A2(n18), .B1(out1[3]), .B2(ci), .ZN(n6) );
  INV_X1 U5 ( .A(n7), .ZN(s[2]) );
  AOI22_X1 U6 ( .A1(out0[2]), .A2(n18), .B1(out1[2]), .B2(ci), .ZN(n7) );
  INV_X1 U7 ( .A(n8), .ZN(s[1]) );
  AOI22_X1 U8 ( .A1(out0[1]), .A2(n18), .B1(out1[1]), .B2(ci), .ZN(n8) );
  INV_X1 U9 ( .A(n9), .ZN(s[0]) );
  AOI22_X1 U10 ( .A1(out0[0]), .A2(n18), .B1(out1[0]), .B2(ci), .ZN(n9) );
  INV_X1 U11 ( .A(ci), .ZN(n18) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_7 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n6, n7, n8, n9, n26;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(n8), .ZN(s[1]) );
  INV_X1 U4 ( .A(n6), .ZN(s[3]) );
  INV_X1 U5 ( .A(n7), .ZN(s[2]) );
  INV_X1 U6 ( .A(n9), .ZN(s[0]) );
  AOI22_X1 U7 ( .A1(out0[1]), .A2(n26), .B1(out1[1]), .B2(ci), .ZN(n8) );
  AOI22_X1 U8 ( .A1(out0[0]), .A2(n26), .B1(out1[0]), .B2(ci), .ZN(n9) );
  AOI22_X1 U9 ( .A1(out0[2]), .A2(n26), .B1(out1[2]), .B2(ci), .ZN(n7) );
  AOI22_X1 U10 ( .A1(out0[3]), .A2(n26), .B1(out1[3]), .B2(ci), .ZN(n6) );
  INV_X1 U11 ( .A(ci), .ZN(n26) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_6 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n26, n27, n28, n29, n30;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(n30), .ZN(s[3]) );
  INV_X1 U4 ( .A(n29), .ZN(s[2]) );
  INV_X1 U5 ( .A(n28), .ZN(s[1]) );
  INV_X1 U6 ( .A(n27), .ZN(s[0]) );
  AOI22_X1 U7 ( .A1(out0[3]), .A2(n26), .B1(out1[3]), .B2(ci), .ZN(n30) );
  AOI22_X1 U8 ( .A1(out0[0]), .A2(n26), .B1(out1[0]), .B2(ci), .ZN(n27) );
  AOI22_X1 U9 ( .A1(out0[1]), .A2(n26), .B1(out1[1]), .B2(ci), .ZN(n28) );
  AOI22_X1 U10 ( .A1(out0[2]), .A2(n26), .B1(out1[2]), .B2(ci), .ZN(n29) );
  INV_X1 U11 ( .A(ci), .ZN(n26) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_5 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n26, n27, n28, n29, n30;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(ci), .ZN(n26) );
  INV_X1 U4 ( .A(n28), .ZN(s[1]) );
  AOI22_X1 U5 ( .A1(out0[1]), .A2(n26), .B1(out1[1]), .B2(ci), .ZN(n28) );
  INV_X1 U6 ( .A(n29), .ZN(s[2]) );
  AOI22_X1 U7 ( .A1(out0[2]), .A2(n26), .B1(out1[2]), .B2(ci), .ZN(n29) );
  INV_X1 U8 ( .A(n30), .ZN(s[3]) );
  AOI22_X1 U9 ( .A1(out0[3]), .A2(n26), .B1(out1[3]), .B2(ci), .ZN(n30) );
  INV_X1 U10 ( .A(n27), .ZN(s[0]) );
  AOI22_X1 U11 ( .A1(out0[0]), .A2(n26), .B1(out1[0]), .B2(ci), .ZN(n27) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_4 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n26, n27, n28, n29, n30;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  INV_X1 U3 ( .A(n30), .ZN(s[3]) );
  INV_X1 U4 ( .A(n29), .ZN(s[2]) );
  INV_X1 U5 ( .A(n28), .ZN(s[1]) );
  INV_X1 U6 ( .A(n27), .ZN(s[0]) );
  AOI22_X1 U7 ( .A1(out0[3]), .A2(n26), .B1(out1[3]), .B2(ci), .ZN(n30) );
  AOI22_X1 U8 ( .A1(out0[2]), .A2(n26), .B1(out1[2]), .B2(ci), .ZN(n29) );
  AOI22_X1 U9 ( .A1(out0[1]), .A2(n26), .B1(out1[1]), .B2(ci), .ZN(n28) );
  AOI22_X1 U10 ( .A1(out0[0]), .A2(n26), .B1(out1[0]), .B2(ci), .ZN(n27) );
  INV_X1 U11 ( .A(ci), .ZN(n26) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_3 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n26, n27, n28, n29;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  MUX2_X1 U3 ( .A(out0[1]), .B(out1[1]), .S(ci), .Z(s[1]) );
  INV_X1 U4 ( .A(n27), .ZN(s[0]) );
  AOI22_X1 U5 ( .A1(out0[3]), .A2(n26), .B1(out1[3]), .B2(ci), .ZN(n29) );
  AOI22_X1 U6 ( .A1(out0[2]), .A2(n26), .B1(out1[2]), .B2(ci), .ZN(n28) );
  AOI22_X1 U7 ( .A1(out0[0]), .A2(n26), .B1(out1[0]), .B2(ci), .ZN(n27) );
  INV_X1 U8 ( .A(ci), .ZN(n26) );
  INV_X1 U9 ( .A(n28), .ZN(s[2]) );
  INV_X1 U10 ( .A(n29), .ZN(s[3]) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_2 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n26, n27, n28, n29, n30;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  AOI22_X1 U3 ( .A1(out0[3]), .A2(n26), .B1(out1[3]), .B2(ci), .ZN(n30) );
  AOI22_X1 U4 ( .A1(out0[2]), .A2(n26), .B1(out1[2]), .B2(ci), .ZN(n29) );
  AOI22_X1 U5 ( .A1(out0[1]), .A2(n26), .B1(out1[1]), .B2(ci), .ZN(n28) );
  AOI22_X1 U6 ( .A1(out0[0]), .A2(n26), .B1(out1[0]), .B2(ci), .ZN(n27) );
  INV_X1 U7 ( .A(ci), .ZN(n26) );
  INV_X1 U8 ( .A(n29), .ZN(s[2]) );
  INV_X1 U9 ( .A(n28), .ZN(s[1]) );
  INV_X1 U10 ( .A(n27), .ZN(s[0]) );
  INV_X1 U11 ( .A(n30), .ZN(s[3]) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12;

  XOR2_X1 U3 ( .A(Ci), .B(n11), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  INV_X1 U1 ( .A(n12), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n11), .B2(Ci), .ZN(n12) );
endmodule


module RCA_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSb_1 ( A, B, ci, s );
  input [3:0] A;
  input [3:0] B;
  output [3:0] s;
  input ci;
  wire   n26, n27, n28, n29, n30;
  wire   [3:0] out0;
  wire   [3:0] out1;

  RCA_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(out0) );
  RCA_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(out1) );
  AOI22_X1 U3 ( .A1(out0[3]), .A2(n26), .B1(out1[3]), .B2(ci), .ZN(n30) );
  AOI22_X1 U4 ( .A1(out0[2]), .A2(n26), .B1(out1[2]), .B2(ci), .ZN(n29) );
  AOI22_X1 U5 ( .A1(out0[1]), .A2(n26), .B1(out1[1]), .B2(ci), .ZN(n28) );
  AOI22_X1 U6 ( .A1(out0[0]), .A2(n26), .B1(out1[0]), .B2(ci), .ZN(n27) );
  INV_X1 U7 ( .A(ci), .ZN(n26) );
  INV_X1 U8 ( .A(n27), .ZN(s[0]) );
  INV_X1 U9 ( .A(n28), .ZN(s[1]) );
  INV_X1 U10 ( .A(n29), .ZN(s[2]) );
  INV_X1 U11 ( .A(n30), .ZN(s[3]) );
endmodule


module CSA ( A, B, c, s );
  input [31:0] A;
  input [31:0] B;
  input [7:0] c;
  output [31:0] s;


  CSb_0 CSbi_0 ( .A(A[3:0]), .B(B[3:0]), .ci(c[0]), .s(s[3:0]) );
  CSb_7 CSbi_1 ( .A(A[7:4]), .B(B[7:4]), .ci(c[1]), .s(s[7:4]) );
  CSb_6 CSbi_2 ( .A(A[11:8]), .B(B[11:8]), .ci(c[2]), .s(s[11:8]) );
  CSb_5 CSbi_3 ( .A(A[15:12]), .B(B[15:12]), .ci(c[3]), .s(s[15:12]) );
  CSb_4 CSbi_4 ( .A(A[19:16]), .B(B[19:16]), .ci(c[4]), .s(s[19:16]) );
  CSb_3 CSbi_5 ( .A(A[23:20]), .B(B[23:20]), .ci(c[5]), .s(s[23:20]) );
  CSb_2 CSbi_6 ( .A(A[27:24]), .B(B[27:24]), .ci(c[6]), .s(s[27:24]) );
  CSb_1 CSbi_7 ( .A(A[31:28]), .B(B[31:28]), .ci(c[7]), .s(s[31:28]) );
endmodule


module P4ADDER_n_bit32 ( A, B, cin0, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input cin0;
  wire   n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;
  wire   [7:1] carries;
  wire   [31:0] BS;
  wire   SYNOPSYS_UNCONNECTED__0;

  XOR2_X1 U3 ( .A(n17), .B(B[8]), .Z(BS[8]) );
  XOR2_X1 U4 ( .A(n17), .B(B[7]), .Z(BS[7]) );
  XOR2_X1 U5 ( .A(n17), .B(B[6]), .Z(BS[6]) );
  XOR2_X1 U6 ( .A(n17), .B(B[5]), .Z(BS[5]) );
  XOR2_X1 U7 ( .A(n17), .B(B[4]), .Z(BS[4]) );
  XOR2_X1 U9 ( .A(n17), .B(B[31]), .Z(BS[31]) );
  XOR2_X1 U10 ( .A(n17), .B(B[30]), .Z(BS[30]) );
  XOR2_X1 U11 ( .A(n17), .B(B[2]), .Z(BS[2]) );
  XOR2_X1 U12 ( .A(n17), .B(B[29]), .Z(BS[29]) );
  XOR2_X1 U13 ( .A(n17), .B(B[28]), .Z(BS[28]) );
  XOR2_X1 U14 ( .A(n17), .B(B[27]), .Z(BS[27]) );
  XOR2_X1 U15 ( .A(n17), .B(B[26]), .Z(BS[26]) );
  XOR2_X1 U16 ( .A(n17), .B(B[25]), .Z(BS[25]) );
  XOR2_X1 U17 ( .A(n17), .B(B[24]), .Z(BS[24]) );
  XOR2_X1 U18 ( .A(n17), .B(B[23]), .Z(BS[23]) );
  XOR2_X1 U19 ( .A(n17), .B(B[22]), .Z(BS[22]) );
  XOR2_X1 U20 ( .A(n17), .B(B[21]), .Z(BS[21]) );
  XOR2_X1 U21 ( .A(n17), .B(B[20]), .Z(BS[20]) );
  XOR2_X1 U22 ( .A(n17), .B(B[1]), .Z(BS[1]) );
  XOR2_X1 U23 ( .A(n17), .B(B[19]), .Z(BS[19]) );
  XOR2_X1 U24 ( .A(n17), .B(B[18]), .Z(BS[18]) );
  XOR2_X1 U25 ( .A(n17), .B(B[17]), .Z(BS[17]) );
  XOR2_X1 U26 ( .A(n17), .B(B[16]), .Z(BS[16]) );
  XOR2_X1 U27 ( .A(n17), .B(B[15]), .Z(BS[15]) );
  XOR2_X1 U28 ( .A(n17), .B(B[14]), .Z(BS[14]) );
  XOR2_X1 U29 ( .A(n17), .B(B[13]), .Z(BS[13]) );
  XOR2_X1 U30 ( .A(n17), .B(B[12]), .Z(BS[12]) );
  XOR2_X1 U31 ( .A(n17), .B(B[11]), .Z(BS[11]) );
  XOR2_X1 U32 ( .A(n17), .B(B[10]), .Z(BS[10]) );
  Cg CG1 ( .A(A), .B({BS[31:1], n1}), .cin0(n17), .cout({
        SYNOPSYS_UNCONNECTED__0, carries}) );
  CSA CSA1 ( .A(A), .B({BS[31:16], n15, n5, n7, BS[12], n14, BS[10], n13, 
        BS[8], n6, BS[6], n4, BS[4], n12, BS[2], n11, n16}), .c({carries, n17}), .s(S) );
  BUF_X4 U1 ( .A(cin0), .Z(n17) );
  CLKBUF_X1 U2 ( .A(BS[5]), .Z(n4) );
  XNOR2_X1 U8 ( .A(n8), .B(B[9]), .ZN(BS[9]) );
  XNOR2_X1 U33 ( .A(n8), .B(B[0]), .ZN(n1) );
  XOR2_X1 U34 ( .A(n17), .B(B[14]), .Z(n5) );
  XOR2_X1 U35 ( .A(n17), .B(B[7]), .Z(n6) );
  XOR2_X1 U36 ( .A(n17), .B(B[13]), .Z(n7) );
  OR2_X1 U37 ( .A1(B[3]), .A2(n8), .ZN(n9) );
  INV_X1 U38 ( .A(cin0), .ZN(n8) );
  NAND2_X1 U39 ( .A1(B[3]), .A2(n8), .ZN(n10) );
  NAND2_X1 U40 ( .A1(n9), .A2(n10), .ZN(BS[3]) );
  CLKBUF_X1 U41 ( .A(BS[1]), .Z(n11) );
  CLKBUF_X1 U42 ( .A(BS[3]), .Z(n12) );
  CLKBUF_X1 U43 ( .A(n1), .Z(n16) );
  BUF_X1 U44 ( .A(BS[9]), .Z(n13) );
  BUF_X1 U45 ( .A(BS[11]), .Z(n14) );
  BUF_X1 U46 ( .A(BS[15]), .Z(n15) );
endmodule


module COMPARATOR_M32_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n26, n27, n29, n30, n31, n32, n33, n34,
         n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n55, n56, n58, n59, n60, n61, n62, n63, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n82, n83,
         n86, n88, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n100,
         n101, n103, n105, n106, n107, n108, n109, n110, n111, n112, n115,
         n116, n118, n119, n120, n121, n122, n123, n124, n125, n126, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n141,
         n142, n144, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n159, n161, n162, n163, n164, n165, n167, n168, n169,
         n172, n175, n176, n177, n178, n179, n180, n181, n182, n183, n193,
         n194, n195, n198, n200, n201, n204, n206, n207, n208, n209, n210,
         n211, n212, n216, n218, n225, n226, n227, n228, n231, n233, n234,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n255, n256,
         n257, n258, n263, n264, n268, n269, n270, n271, n272, n273, n276,
         n278, n286, n287, n288, n289, n290, n292, n293, n294, n295, n298,
         n300, n301, n303, n305, n306, n313, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511;

  NAND3_X1 U281 ( .A1(n16), .A2(n17), .A3(n15), .ZN(n11) );
  NAND3_X1 U282 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n20) );
  NAND3_X1 U283 ( .A1(n425), .A2(n29), .A3(n418), .ZN(n22) );
  NAND3_X1 U284 ( .A1(n39), .A2(n429), .A3(n40), .ZN(n43) );
  NAND3_X1 U285 ( .A1(n40), .A2(n52), .A3(n53), .ZN(n51) );
  NAND3_X1 U286 ( .A1(n438), .A2(n58), .A3(n432), .ZN(n52) );
  NAND3_X1 U287 ( .A1(n60), .A2(n39), .A3(n61), .ZN(n50) );
  NAND3_X1 U288 ( .A1(n76), .A2(n77), .A3(n78), .ZN(n75) );
  NAND3_X1 U289 ( .A1(n97), .A2(n457), .A3(n98), .ZN(n101) );
  NAND3_X1 U292 ( .A1(n467), .A2(n460), .A3(n118), .ZN(n111) );
  NAND3_X1 U293 ( .A1(n120), .A2(n97), .A3(n121), .ZN(n109) );
  NAND3_X1 U294 ( .A1(n132), .A2(n137), .A3(n138), .ZN(n123) );
  NAND3_X1 U295 ( .A1(n478), .A2(n144), .A3(n473), .ZN(n137) );
  NAND3_X1 U296 ( .A1(n151), .A2(n152), .A3(n153), .ZN(n147) );
  NAND3_X1 U297 ( .A1(n167), .A2(n168), .A3(n169), .ZN(n164) );
  NAND3_X1 U298 ( .A1(n27), .A2(n418), .A3(n423), .ZN(n167) );
  NAND3_X1 U299 ( .A1(n183), .A2(n431), .A3(n46), .ZN(n182) );
  NAND3_X1 U300 ( .A1(n183), .A2(n46), .A3(n41), .ZN(n180) );
  NAND3_X1 U301 ( .A1(n436), .A2(n56), .A3(n432), .ZN(n195) );
  NAND3_X1 U304 ( .A1(n216), .A2(n70), .A3(n72), .ZN(n211) );
  NAND3_X1 U305 ( .A1(n218), .A2(n1), .A3(n432), .ZN(n209) );
  NAND3_X1 U307 ( .A1(n216), .A2(n444), .A3(n70), .ZN(n218) );
  NAND3_X1 U308 ( .A1(n245), .A2(n459), .A3(n105), .ZN(n244) );
  NAND3_X1 U309 ( .A1(n245), .A2(n105), .A3(n99), .ZN(n242) );
  NAND3_X1 U310 ( .A1(n464), .A2(n116), .A3(n460), .ZN(n257) );
  NAND3_X1 U311 ( .A1(n276), .A2(n136), .A3(n133), .ZN(n272) );
  NAND3_X1 U312 ( .A1(n278), .A2(n465), .A3(n460), .ZN(n270) );
  NAND3_X1 U313 ( .A1(n276), .A2(n472), .A3(n136), .ZN(n278) );
  NAND3_X1 U314 ( .A1(n286), .A2(n287), .A3(n288), .ZN(n268) );
  NAND3_X1 U315 ( .A1(n293), .A2(n294), .A3(n295), .ZN(n287) );
  AOI21_X1 U1 ( .B1(n176), .B2(n177), .A(n178), .ZN(n163) );
  NAND4_X1 U2 ( .A1(n179), .A2(n180), .A3(n181), .A4(n182), .ZN(n178) );
  AND3_X1 U3 ( .A1(n193), .A2(n194), .A3(n195), .ZN(n177) );
  OAI21_X1 U4 ( .B1(n206), .B2(n207), .A(n208), .ZN(n176) );
  AOI21_X1 U5 ( .B1(n238), .B2(n239), .A(n240), .ZN(n206) );
  NAND4_X1 U6 ( .A1(n241), .A2(n242), .A3(n243), .A4(n244), .ZN(n240) );
  NAND2_X1 U7 ( .A1(n268), .A2(n269), .ZN(n238) );
  NOR2_X1 U8 ( .A1(n255), .A2(n256), .ZN(n239) );
  OAI21_X1 U9 ( .B1(n47), .B2(n48), .A(n49), .ZN(n18) );
  NAND2_X1 U10 ( .A1(n62), .A2(n63), .ZN(n48) );
  NOR2_X1 U11 ( .A1(n50), .A2(n51), .ZN(n49) );
  AOI21_X1 U12 ( .B1(n73), .B2(n74), .A(n75), .ZN(n47) );
  INV_X1 U13 ( .A(n55), .ZN(n432) );
  NOR2_X1 U14 ( .A1(n96), .A2(n83), .ZN(n243) );
  NOR2_X1 U15 ( .A1(n38), .A2(n26), .ZN(n181) );
  NOR2_X1 U16 ( .A1(n83), .A2(n448), .ZN(n79) );
  INV_X1 U17 ( .A(n26), .ZN(n418) );
  NOR2_X1 U18 ( .A1(n96), .A2(n83), .ZN(n95) );
  NOR2_X1 U19 ( .A1(n209), .A2(n210), .ZN(n208) );
  NAND2_X1 U20 ( .A1(n211), .A2(n212), .ZN(n210) );
  NOR2_X1 U21 ( .A1(n441), .A2(n435), .ZN(n212) );
  NOR2_X1 U22 ( .A1(n38), .A2(n26), .ZN(n37) );
  NOR2_X1 U23 ( .A1(n130), .A2(n115), .ZN(n129) );
  NOR2_X1 U24 ( .A1(n447), .A2(n88), .ZN(n76) );
  NAND2_X1 U25 ( .A1(n450), .A2(n445), .ZN(n77) );
  AOI21_X1 U26 ( .B1(n79), .B2(n452), .A(n441), .ZN(n78) );
  INV_X1 U27 ( .A(n115), .ZN(n460) );
  NOR2_X1 U28 ( .A1(n141), .A2(n154), .ZN(n153) );
  NOR2_X1 U29 ( .A1(n141), .A2(n154), .ZN(n295) );
  INV_X1 U30 ( .A(n83), .ZN(n445) );
  INV_X1 U31 ( .A(n141), .ZN(n473) );
  INV_X1 U32 ( .A(n8), .ZN(LE) );
  INV_X1 U33 ( .A(n99), .ZN(n455) );
  INV_X1 U34 ( .A(n133), .ZN(n469) );
  INV_X1 U35 ( .A(n41), .ZN(n427) );
  INV_X1 U36 ( .A(n130), .ZN(n465) );
  OAI21_X1 U37 ( .B1(n10), .B2(n11), .A(n12), .ZN(n8) );
  NOR2_X1 U38 ( .A1(n13), .A2(n3), .ZN(n12) );
  AOI21_X1 U39 ( .B1(n18), .B2(n19), .A(n20), .ZN(n10) );
  NAND2_X1 U40 ( .A1(n90), .A2(n231), .ZN(n83) );
  NAND2_X1 U41 ( .A1(n150), .A2(n298), .ZN(n141) );
  INV_X1 U42 ( .A(n120), .ZN(n459) );
  INV_X1 U43 ( .A(n60), .ZN(n431) );
  NAND4_X1 U44 ( .A1(n105), .A2(n103), .A3(n245), .A4(n264), .ZN(n255) );
  NAND2_X1 U45 ( .A1(n32), .A2(n172), .ZN(n26) );
  INV_X1 U46 ( .A(n45), .ZN(n429) );
  NAND2_X1 U47 ( .A1(n121), .A2(n264), .ZN(n115) );
  NOR2_X1 U48 ( .A1(n270), .A2(n271), .ZN(n269) );
  NAND2_X1 U49 ( .A1(n272), .A2(n273), .ZN(n271) );
  NOR2_X1 U50 ( .A1(n83), .A2(n106), .ZN(n234) );
  NOR2_X1 U51 ( .A1(n91), .A2(n92), .ZN(n74) );
  NAND2_X1 U52 ( .A1(n100), .A2(n101), .ZN(n91) );
  OAI21_X1 U53 ( .B1(n455), .B2(n94), .A(n95), .ZN(n92) );
  NOR2_X1 U54 ( .A1(n33), .A2(n34), .ZN(n19) );
  NAND2_X1 U55 ( .A1(n42), .A2(n43), .ZN(n33) );
  OAI21_X1 U56 ( .B1(n427), .B2(n36), .A(n37), .ZN(n34) );
  AND2_X1 U57 ( .A1(n29), .A2(n46), .ZN(n42) );
  NOR2_X1 U58 ( .A1(n141), .A2(n144), .ZN(n290) );
  NOR2_X1 U59 ( .A1(n439), .A2(n65), .ZN(n63) );
  INV_X1 U60 ( .A(n70), .ZN(n439) );
  OAI21_X1 U61 ( .B1(n66), .B2(n67), .A(n58), .ZN(n65) );
  NAND2_X1 U62 ( .A1(n68), .A2(n69), .ZN(n67) );
  NOR2_X1 U63 ( .A1(n141), .A2(n292), .ZN(n289) );
  NAND2_X1 U64 ( .A1(n435), .A2(n432), .ZN(n53) );
  INV_X1 U65 ( .A(n59), .ZN(n438) );
  AND2_X1 U66 ( .A1(n16), .A2(n172), .ZN(n168) );
  NAND2_X1 U67 ( .A1(n420), .A2(n418), .ZN(n169) );
  NAND2_X1 U68 ( .A1(n476), .A2(n473), .ZN(n138) );
  INV_X1 U69 ( .A(n146), .ZN(n478) );
  NOR2_X1 U70 ( .A1(n125), .A2(n126), .ZN(n124) );
  OAI211_X1 U71 ( .C1(n134), .C2(n135), .A(n118), .B(n136), .ZN(n125) );
  OAI21_X1 U72 ( .B1(n469), .B2(n128), .A(n129), .ZN(n126) );
  NAND2_X1 U73 ( .A1(n132), .A2(n131), .ZN(n135) );
  NOR2_X1 U74 ( .A1(n450), .A2(n237), .ZN(n233) );
  AND2_X1 U75 ( .A1(n31), .A2(n32), .ZN(n21) );
  NAND2_X1 U76 ( .A1(n422), .A2(n418), .ZN(n23) );
  NOR2_X1 U77 ( .A1(n448), .A2(n453), .ZN(n100) );
  INV_X1 U78 ( .A(n105), .ZN(n453) );
  NOR2_X1 U79 ( .A1(n2), .A2(n71), .ZN(n62) );
  AND3_X1 U80 ( .A1(n69), .A2(n68), .A3(n72), .ZN(n2) );
  NAND2_X1 U81 ( .A1(n432), .A2(n1), .ZN(n71) );
  NOR2_X1 U82 ( .A1(n305), .A2(n306), .ZN(n286) );
  AOI21_X1 U83 ( .B1(n289), .B2(n142), .A(n290), .ZN(n288) );
  INV_X1 U84 ( .A(n89), .ZN(n444) );
  NAND2_X1 U85 ( .A1(n39), .A2(n183), .ZN(n41) );
  NAND2_X1 U86 ( .A1(n146), .A2(n292), .ZN(n154) );
  NAND2_X1 U87 ( .A1(n97), .A2(n245), .ZN(n99) );
  NAND2_X1 U88 ( .A1(n82), .A2(n237), .ZN(n96) );
  NOR2_X1 U89 ( .A1(n9), .A2(n8), .ZN(EQ) );
  NAND2_X1 U90 ( .A1(n131), .A2(n276), .ZN(n133) );
  NAND2_X1 U91 ( .A1(n30), .A2(n175), .ZN(n38) );
  NAND2_X1 U92 ( .A1(n119), .A2(n263), .ZN(n130) );
  NAND2_X1 U93 ( .A1(n61), .A2(n204), .ZN(n55) );
  INV_X1 U94 ( .A(n68), .ZN(n441) );
  NAND2_X1 U95 ( .A1(n69), .A2(n216), .ZN(n72) );
  NAND2_X1 U96 ( .A1(n89), .A2(n69), .ZN(n88) );
  INV_X1 U97 ( .A(n198), .ZN(n436) );
  NOR2_X1 U98 ( .A1(n200), .A2(n201), .ZN(n193) );
  NAND2_X1 U99 ( .A1(n183), .A2(n204), .ZN(n200) );
  NAND2_X1 U100 ( .A1(n46), .A2(n45), .ZN(n201) );
  NAND2_X1 U101 ( .A1(n70), .A2(n66), .ZN(n228) );
  INV_X1 U102 ( .A(n56), .ZN(n435) );
  INV_X1 U103 ( .A(n86), .ZN(n450) );
  NAND2_X1 U104 ( .A1(n131), .A2(n132), .ZN(n128) );
  INV_X1 U105 ( .A(n106), .ZN(n448) );
  NAND2_X1 U106 ( .A1(n39), .A2(n40), .ZN(n36) );
  NAND2_X1 U107 ( .A1(n97), .A2(n98), .ZN(n94) );
  NAND2_X1 U108 ( .A1(n276), .A2(n298), .ZN(n305) );
  NAND2_X1 U109 ( .A1(n136), .A2(n134), .ZN(n306) );
  AND2_X1 U110 ( .A1(n59), .A2(n198), .ZN(n1) );
  INV_X1 U111 ( .A(n82), .ZN(n452) );
  NAND2_X1 U112 ( .A1(n257), .A2(n258), .ZN(n256) );
  NAND2_X1 U113 ( .A1(n462), .A2(n460), .ZN(n258) );
  INV_X1 U114 ( .A(n263), .ZN(n464) );
  NAND2_X1 U115 ( .A1(n111), .A2(n112), .ZN(n110) );
  AND2_X1 U116 ( .A1(n313), .A2(n98), .ZN(n112) );
  OR2_X1 U117 ( .A1(n115), .A2(n116), .ZN(n313) );
  NAND2_X1 U118 ( .A1(n225), .A2(n226), .ZN(n207) );
  NOR2_X1 U119 ( .A1(n227), .A2(n228), .ZN(n226) );
  AOI21_X1 U120 ( .B1(n233), .B2(n445), .A(n234), .ZN(n225) );
  NAND2_X1 U121 ( .A1(n216), .A2(n231), .ZN(n227) );
  INV_X1 U122 ( .A(n27), .ZN(n422) );
  INV_X1 U123 ( .A(n118), .ZN(n462) );
  INV_X1 U124 ( .A(n90), .ZN(n447) );
  INV_X1 U125 ( .A(n142), .ZN(n476) );
  NAND2_X1 U126 ( .A1(n107), .A2(n108), .ZN(n73) );
  NOR2_X1 U127 ( .A1(n109), .A2(n110), .ZN(n108) );
  OAI21_X1 U128 ( .B1(n122), .B2(n123), .A(n124), .ZN(n107) );
  NAND2_X1 U129 ( .A1(n147), .A2(n148), .ZN(n122) );
  AND2_X1 U130 ( .A1(n150), .A2(n6), .ZN(n148) );
  AND2_X1 U131 ( .A1(n149), .A2(n131), .ZN(n6) );
  AND2_X1 U132 ( .A1(n5), .A2(n15), .ZN(n165) );
  AND2_X1 U133 ( .A1(n31), .A2(n17), .ZN(n5) );
  AND2_X1 U134 ( .A1(n132), .A2(n116), .ZN(n273) );
  AND2_X1 U135 ( .A1(n40), .A2(n27), .ZN(n179) );
  AND2_X1 U136 ( .A1(n98), .A2(n86), .ZN(n241) );
  INV_X1 U137 ( .A(n30), .ZN(n425) );
  INV_X1 U138 ( .A(n119), .ZN(n467) );
  INV_X1 U139 ( .A(n29), .ZN(n420) );
  OR2_X1 U140 ( .A1(n58), .A2(n55), .ZN(n194) );
  INV_X1 U141 ( .A(n149), .ZN(n472) );
  INV_X1 U142 ( .A(n9), .ZN(GE) );
  INV_X1 U143 ( .A(n103), .ZN(n457) );
  INV_X1 U144 ( .A(n175), .ZN(n423) );
  INV_X1 U145 ( .A(A[6]), .ZN(n470) );
  INV_X1 U146 ( .A(A[24]), .ZN(n428) );
  INV_X1 U147 ( .A(A[25]), .ZN(n426) );
  NAND2_X1 U148 ( .A1(A[18]), .A2(n493), .ZN(n69) );
  NAND2_X1 U149 ( .A1(A[6]), .A2(n505), .ZN(n131) );
  NAND2_X1 U150 ( .A1(A[7]), .A2(n504), .ZN(n132) );
  NAND2_X1 U151 ( .A1(A[12]), .A2(n499), .ZN(n97) );
  NAND2_X1 U152 ( .A1(A[24]), .A2(n487), .ZN(n39) );
  NAND2_X1 U153 ( .A1(A[25]), .A2(n486), .ZN(n40) );
  INV_X1 U154 ( .A(A[21]), .ZN(n434) );
  NAND2_X1 U155 ( .A1(A[13]), .A2(n498), .ZN(n98) );
  INV_X1 U156 ( .A(A[22]), .ZN(n433) );
  INV_X1 U157 ( .A(B[2]), .ZN(n509) );
  INV_X1 U158 ( .A(A[14]), .ZN(n451) );
  INV_X1 U159 ( .A(A[23]), .ZN(n430) );
  NAND2_X1 U160 ( .A1(A[19]), .A2(n492), .ZN(n68) );
  NAND2_X1 U161 ( .A1(A[27]), .A2(n484), .ZN(n27) );
  INV_X1 U162 ( .A(B[27]), .ZN(n484) );
  NAND2_X1 U163 ( .A1(A[3]), .A2(n508), .ZN(n142) );
  INV_X1 U164 ( .A(B[3]), .ZN(n508) );
  NAND2_X1 U165 ( .A1(A[26]), .A2(n485), .ZN(n30) );
  INV_X1 U166 ( .A(B[26]), .ZN(n485) );
  NAND2_X1 U167 ( .A1(A[8]), .A2(n503), .ZN(n119) );
  INV_X1 U168 ( .A(B[8]), .ZN(n503) );
  NAND2_X1 U169 ( .A1(A[14]), .A2(n497), .ZN(n82) );
  NAND2_X1 U170 ( .A1(A[17]), .A2(n494), .ZN(n89) );
  INV_X1 U171 ( .A(B[17]), .ZN(n494) );
  INV_X1 U172 ( .A(B[4]), .ZN(n507) );
  NAND2_X1 U173 ( .A1(A[16]), .A2(n495), .ZN(n90) );
  INV_X1 U174 ( .A(A[28]), .ZN(n419) );
  NAND2_X1 U175 ( .A1(A[23]), .A2(n488), .ZN(n60) );
  NAND2_X1 U176 ( .A1(A[9]), .A2(n502), .ZN(n116) );
  NAND2_X1 U177 ( .A1(A[22]), .A2(n489), .ZN(n61) );
  NAND2_X1 U178 ( .A1(n161), .A2(n162), .ZN(n9) );
  NOR2_X1 U179 ( .A1(n4), .A2(n7), .ZN(n161) );
  OAI21_X1 U180 ( .B1(n163), .B2(n164), .A(n165), .ZN(n162) );
  NAND2_X1 U181 ( .A1(A[15]), .A2(n496), .ZN(n86) );
  NAND2_X1 U182 ( .A1(A[21]), .A2(n490), .ZN(n56) );
  NAND2_X1 U183 ( .A1(A[28]), .A2(n483), .ZN(n32) );
  NAND2_X1 U184 ( .A1(A[11]), .A2(n500), .ZN(n120) );
  NAND2_X1 U185 ( .A1(A[20]), .A2(n491), .ZN(n59) );
  NAND2_X1 U186 ( .A1(A[5]), .A2(n506), .ZN(n149) );
  INV_X1 U187 ( .A(B[5]), .ZN(n506) );
  NAND2_X1 U188 ( .A1(A[29]), .A2(n482), .ZN(n31) );
  INV_X1 U189 ( .A(A[1]), .ZN(n479) );
  INV_X1 U190 ( .A(A[30]), .ZN(n416) );
  INV_X1 U191 ( .A(A[29]), .ZN(n417) );
  NAND2_X1 U192 ( .A1(B[27]), .A2(n421), .ZN(n29) );
  INV_X1 U193 ( .A(A[27]), .ZN(n421) );
  NAND2_X1 U194 ( .A1(B[4]), .A2(n474), .ZN(n298) );
  NAND2_X1 U195 ( .A1(B[2]), .A2(n477), .ZN(n292) );
  NAND2_X1 U196 ( .A1(B[26]), .A2(n424), .ZN(n175) );
  INV_X1 U197 ( .A(A[26]), .ZN(n424) );
  NAND2_X1 U198 ( .A1(B[17]), .A2(n443), .ZN(n66) );
  INV_X1 U199 ( .A(A[17]), .ZN(n443) );
  NAND2_X1 U200 ( .A1(B[8]), .A2(n466), .ZN(n263) );
  INV_X1 U201 ( .A(A[8]), .ZN(n466) );
  NAND2_X1 U202 ( .A1(B[5]), .A2(n471), .ZN(n134) );
  INV_X1 U203 ( .A(A[5]), .ZN(n471) );
  INV_X1 U204 ( .A(A[31]), .ZN(n415) );
  NAND2_X1 U205 ( .A1(B[3]), .A2(n475), .ZN(n144) );
  INV_X1 U206 ( .A(A[3]), .ZN(n475) );
  INV_X1 U207 ( .A(A[13]), .ZN(n454) );
  INV_X1 U208 ( .A(A[18]), .ZN(n442) );
  INV_X1 U209 ( .A(A[15]), .ZN(n449) );
  INV_X1 U210 ( .A(A[12]), .ZN(n456) );
  INV_X1 U211 ( .A(A[7]), .ZN(n468) );
  INV_X1 U212 ( .A(A[19]), .ZN(n440) );
  INV_X1 U213 ( .A(A[9]), .ZN(n463) );
  INV_X1 U214 ( .A(A[11]), .ZN(n458) );
  INV_X1 U215 ( .A(B[1]), .ZN(n510) );
  AND3_X1 U216 ( .A1(A[30]), .A2(n481), .A3(n15), .ZN(n3) );
  INV_X1 U217 ( .A(A[16]), .ZN(n446) );
  INV_X1 U218 ( .A(A[20]), .ZN(n437) );
  NAND2_X1 U219 ( .A1(n155), .A2(n156), .ZN(n152) );
  NAND2_X1 U220 ( .A1(A[0]), .A2(n511), .ZN(n156) );
  NAND2_X1 U221 ( .A1(A[1]), .A2(n510), .ZN(n155) );
  NAND2_X1 U222 ( .A1(n300), .A2(n301), .ZN(n294) );
  NAND2_X1 U223 ( .A1(B[1]), .A2(n479), .ZN(n300) );
  INV_X1 U224 ( .A(A[0]), .ZN(n480) );
  AND2_X1 U225 ( .A1(n303), .A2(n142), .ZN(n293) );
  NAND2_X1 U226 ( .A1(A[1]), .A2(n510), .ZN(n303) );
  AND2_X1 U227 ( .A1(n159), .A2(n144), .ZN(n151) );
  NAND2_X1 U228 ( .A1(B[1]), .A2(n479), .ZN(n159) );
  NAND2_X1 U229 ( .A1(A[2]), .A2(n509), .ZN(n146) );
  INV_X1 U230 ( .A(A[2]), .ZN(n477) );
  NAND2_X1 U231 ( .A1(A[4]), .A2(n507), .ZN(n150) );
  INV_X1 U232 ( .A(A[4]), .ZN(n474) );
  NAND2_X1 U233 ( .A1(A[10]), .A2(n501), .ZN(n121) );
  INV_X1 U234 ( .A(A[10]), .ZN(n461) );
  NAND2_X1 U235 ( .A1(B[14]), .A2(n451), .ZN(n237) );
  INV_X1 U236 ( .A(B[14]), .ZN(n497) );
  NAND2_X1 U237 ( .A1(B[13]), .A2(n454), .ZN(n105) );
  INV_X1 U238 ( .A(B[13]), .ZN(n498) );
  NAND2_X1 U239 ( .A1(B[12]), .A2(n456), .ZN(n245) );
  INV_X1 U240 ( .A(B[12]), .ZN(n499) );
  AND3_X1 U241 ( .A1(B[30]), .A2(n416), .A3(n15), .ZN(n7) );
  INV_X1 U242 ( .A(B[30]), .ZN(n481) );
  XNOR2_X1 U243 ( .A(B[30]), .B(A[30]), .ZN(n17) );
  NAND2_X1 U244 ( .A1(B[29]), .A2(n417), .ZN(n16) );
  INV_X1 U245 ( .A(B[29]), .ZN(n482) );
  NAND2_X1 U246 ( .A1(B[18]), .A2(n442), .ZN(n216) );
  INV_X1 U247 ( .A(B[18]), .ZN(n493) );
  NAND2_X1 U248 ( .A1(B[9]), .A2(n463), .ZN(n118) );
  INV_X1 U249 ( .A(B[9]), .ZN(n502) );
  NAND2_X1 U250 ( .A1(B[19]), .A2(n440), .ZN(n70) );
  INV_X1 U251 ( .A(B[19]), .ZN(n492) );
  AND2_X1 U252 ( .A1(B[31]), .A2(n415), .ZN(n4) );
  NOR2_X1 U253 ( .A1(B[31]), .A2(n415), .ZN(n13) );
  XNOR2_X1 U254 ( .A(B[31]), .B(A[31]), .ZN(n15) );
  NAND2_X1 U255 ( .A1(B[7]), .A2(n468), .ZN(n136) );
  INV_X1 U256 ( .A(B[7]), .ZN(n504) );
  NAND2_X1 U257 ( .A1(B[21]), .A2(n434), .ZN(n58) );
  INV_X1 U258 ( .A(B[21]), .ZN(n490) );
  NAND2_X1 U259 ( .A1(B[15]), .A2(n449), .ZN(n106) );
  INV_X1 U260 ( .A(B[15]), .ZN(n496) );
  NAND2_X1 U261 ( .A1(B[0]), .A2(n480), .ZN(n301) );
  INV_X1 U262 ( .A(B[0]), .ZN(n511) );
  NAND2_X1 U263 ( .A1(B[16]), .A2(n446), .ZN(n231) );
  INV_X1 U264 ( .A(B[16]), .ZN(n495) );
  NAND2_X1 U265 ( .A1(B[20]), .A2(n437), .ZN(n198) );
  INV_X1 U266 ( .A(B[20]), .ZN(n491) );
  INV_X1 U267 ( .A(B[25]), .ZN(n486) );
  NAND2_X1 U268 ( .A1(B[25]), .A2(n426), .ZN(n46) );
  NAND2_X1 U269 ( .A1(B[11]), .A2(n458), .ZN(n103) );
  INV_X1 U270 ( .A(B[11]), .ZN(n500) );
  NAND2_X1 U271 ( .A1(B[23]), .A2(n430), .ZN(n45) );
  INV_X1 U272 ( .A(B[23]), .ZN(n488) );
  NAND2_X1 U273 ( .A1(B[24]), .A2(n428), .ZN(n183) );
  INV_X1 U274 ( .A(B[24]), .ZN(n487) );
  NAND2_X1 U275 ( .A1(B[10]), .A2(n461), .ZN(n264) );
  INV_X1 U276 ( .A(B[10]), .ZN(n501) );
  NAND2_X1 U277 ( .A1(B[6]), .A2(n470), .ZN(n276) );
  INV_X1 U278 ( .A(B[6]), .ZN(n505) );
  NAND2_X1 U279 ( .A1(B[28]), .A2(n419), .ZN(n172) );
  INV_X1 U280 ( .A(B[28]), .ZN(n483) );
  NAND2_X1 U290 ( .A1(B[22]), .A2(n433), .ZN(n204) );
  INV_X1 U291 ( .A(B[22]), .ZN(n489) );
endmodule


module COMPARATOR_M32 ( A, B, sel, OUTPUT );
  input [31:0] A;
  input [31:0] B;
  input [1:0] sel;
  output [31:0] OUTPUT;
  wire   N12, N15, N16, n5, n6, n8, n9;
  assign OUTPUT[1] = 1'b0;
  assign OUTPUT[2] = 1'b0;
  assign OUTPUT[3] = 1'b0;
  assign OUTPUT[4] = 1'b0;
  assign OUTPUT[5] = 1'b0;
  assign OUTPUT[6] = 1'b0;
  assign OUTPUT[7] = 1'b0;
  assign OUTPUT[8] = 1'b0;
  assign OUTPUT[9] = 1'b0;
  assign OUTPUT[10] = 1'b0;
  assign OUTPUT[11] = 1'b0;
  assign OUTPUT[12] = 1'b0;
  assign OUTPUT[13] = 1'b0;
  assign OUTPUT[14] = 1'b0;
  assign OUTPUT[15] = 1'b0;
  assign OUTPUT[16] = 1'b0;
  assign OUTPUT[17] = 1'b0;
  assign OUTPUT[18] = 1'b0;
  assign OUTPUT[19] = 1'b0;
  assign OUTPUT[20] = 1'b0;
  assign OUTPUT[21] = 1'b0;
  assign OUTPUT[22] = 1'b0;
  assign OUTPUT[23] = 1'b0;
  assign OUTPUT[24] = 1'b0;
  assign OUTPUT[25] = 1'b0;
  assign OUTPUT[26] = 1'b0;
  assign OUTPUT[27] = 1'b0;
  assign OUTPUT[28] = 1'b0;
  assign OUTPUT[29] = 1'b0;
  assign OUTPUT[30] = 1'b0;
  assign OUTPUT[31] = 1'b0;

  XOR2_X1 U8 ( .A(n8), .B(N12), .Z(n6) );
  COMPARATOR_M32_DW01_cmp6_1 r61 ( .A(A), .B(B), .TC(1'b0), .EQ(N12), .LE(N16), 
        .GE(N15) );
  INV_X1 U2 ( .A(sel[1]), .ZN(n9) );
  AOI22_X1 U4 ( .A1(N15), .A2(n8), .B1(N16), .B2(sel[0]), .ZN(n5) );
  INV_X1 U5 ( .A(sel[0]), .ZN(n8) );
  OAI22_X1 U6 ( .A1(n5), .A2(n9), .B1(sel[1]), .B2(n6), .ZN(OUTPUT[0]) );
endmodule


module ALU_M32_C4 ( CODE, DATA1, DATA2, OUTALU );
  input [3:0] CODE;
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTALU;
  wire   \Comparison[1] , \COMPARATORout[0] , n70, n71, n72, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n169, n170, n171, n172, net131848,
         net133061, net134759, net134757, net134755, net134765, net134763,
         net134761, net134777, net134775, net134773, net134771, net134769,
         net134767, net134783, net134781, net134779, net134795, net134793,
         net134791, net134789, net134787, net134785, net131887, net131855, n91,
         n90, net131849, n92, n74, n73, n176, n175, n174, n173, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n657, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804;
  wire   [31:0] SHIFTERout;
  wire   [31:0] ADDERout;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  SHIFTER_M32_N5 SHIFTOP ( .A(DATA1), .B({DATA2[31:4], n645, n663, DATA2[1], 
        n685}), .LEFT_RIGHT(CODE[0]), .OUTPUT(SHIFTERout) );
  P4ADDER_n_bit32 ADDSUBOP ( .A(DATA1), .B({DATA2[31], n695, n698, n701, n686, 
        n697, n703, n702, n705, n736, n694, n688, n691, n708, n711, n707, n699, 
        n693, n704, n700, n689, n706, n692, n687, n690, n696, DATA2[5:0]}), 
        .cin0(net133061), .S(ADDERout) );
  COMPARATOR_M32 COMPOP ( .A(DATA1), .B({DATA2[31], n695, n698, n701, n686, 
        n697, n703, n702, n705, n736, n694, n688, n691, n708, n711, n707, n699, 
        n693, n704, n700, n689, n706, n692, n687, n690, n696, DATA2[5:1], n685}), .sel({\Comparison[1] , net131848}), .OUTPUT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, \COMPARATORout[0] }) );
  XOR2_X1 U209 ( .A(CODE[1]), .B(CODE[0]), .Z(n176) );
  INV_X1 U2 ( .A(n801), .ZN(n645) );
  AOI221_X1 U3 ( .B1(net134767), .B2(n744), .C1(DATA1[30]), .C2(net134781), 
        .A(net134785), .ZN(n100) );
  AOI221_X1 U4 ( .B1(net134771), .B2(n762), .C1(DATA1[12]), .C2(net134779), 
        .A(net134789), .ZN(n160) );
  AOI221_X1 U5 ( .B1(net134767), .B2(n767), .C1(DATA1[7]), .C2(net134783), .A(
        net134785), .ZN(n82) );
  AOI221_X1 U6 ( .B1(net134769), .B2(n753), .C1(DATA1[21]), .C2(net134781), 
        .A(net134787), .ZN(n130) );
  AOI221_X1 U7 ( .B1(net134769), .B2(n750), .C1(DATA1[24]), .C2(net134781), 
        .A(net134787), .ZN(n121) );
  AOI221_X1 U8 ( .B1(net134769), .B2(n748), .C1(DATA1[26]), .C2(net134781), 
        .A(net134787), .ZN(n115) );
  AOI221_X1 U9 ( .B1(net134767), .B2(n747), .C1(DATA1[27]), .C2(net134781), 
        .A(net134785), .ZN(n112) );
  INV_X1 U10 ( .A(CODE[0]), .ZN(net133061) );
  NOR2_X1 U11 ( .A1(n90), .A2(net131887), .ZN(n646) );
  NOR2_X1 U12 ( .A1(n91), .A2(net131855), .ZN(n647) );
  AND2_X1 U13 ( .A1(n726), .A2(n725), .ZN(n648) );
  AND2_X1 U14 ( .A1(n728), .A2(n727), .ZN(n649) );
  AND2_X1 U15 ( .A1(n730), .A2(n729), .ZN(n650) );
  AND2_X1 U16 ( .A1(n714), .A2(n713), .ZN(n651) );
  AND2_X1 U17 ( .A1(n742), .A2(n741), .ZN(n652) );
  NOR3_X1 U18 ( .A1(net131848), .A2(CODE[0]), .A3(n174), .ZN(n77) );
  NOR2_X1 U19 ( .A1(n130), .A2(n784), .ZN(n653) );
  NOR2_X1 U20 ( .A1(n129), .A2(n753), .ZN(n654) );
  NOR2_X1 U21 ( .A1(n653), .A2(n654), .ZN(n655) );
  NAND2_X1 U22 ( .A1(n131), .A2(n655), .ZN(OUTALU[21]) );
  BUF_X1 U23 ( .A(DATA2[7]), .Z(n690) );
  BUF_X1 U24 ( .A(DATA2[13]), .Z(n704) );
  NOR2_X1 U25 ( .A1(n646), .A2(n647), .ZN(n657) );
  NAND2_X1 U26 ( .A1(n92), .A2(n657), .ZN(OUTALU[4]) );
  OAI221_X1 U27 ( .B1(n659), .B2(n660), .C1(n661), .C2(n662), .A(n652), .ZN(
        OUTALU[5]) );
  INV_X1 U28 ( .A(SHIFTERout[5]), .ZN(n659) );
  INV_X1 U29 ( .A(n73), .ZN(n660) );
  INV_X1 U30 ( .A(ADDERout[5]), .ZN(n661) );
  INV_X1 U31 ( .A(n74), .ZN(n662) );
  AOI22_X1 U32 ( .A1(SHIFTERout[21]), .A2(n73), .B1(ADDERout[21]), .B2(n74), 
        .ZN(n131) );
  AOI22_X1 U33 ( .A1(SHIFTERout[3]), .A2(n73), .B1(ADDERout[3]), .B2(n74), 
        .ZN(n95) );
  AOI22_X1 U34 ( .A1(SHIFTERout[8]), .A2(n73), .B1(ADDERout[8]), .B2(n74), 
        .ZN(n80) );
  AOI22_X1 U35 ( .A1(SHIFTERout[4]), .A2(n73), .B1(ADDERout[4]), .B2(n74), 
        .ZN(n92) );
  AOI22_X1 U36 ( .A1(SHIFTERout[1]), .A2(n73), .B1(ADDERout[1]), .B2(n74), 
        .ZN(n137) );
  NAND2_X1 U37 ( .A1(n128), .A2(n648), .ZN(OUTALU[22]) );
  CLKBUF_X1 U38 ( .A(DATA2[2]), .Z(n663) );
  OR2_X1 U39 ( .A1(n120), .A2(n750), .ZN(n664) );
  OR2_X1 U40 ( .A1(n121), .A2(n781), .ZN(n665) );
  NAND3_X1 U41 ( .A1(n664), .A2(n665), .A3(n122), .ZN(OUTALU[24]) );
  BUF_X1 U42 ( .A(DATA2[15]), .Z(n699) );
  OR2_X1 U43 ( .A1(n96), .A2(n743), .ZN(n666) );
  OR2_X1 U44 ( .A1(n97), .A2(n774), .ZN(n667) );
  NAND3_X1 U45 ( .A1(n98), .A2(n667), .A3(n666), .ZN(OUTALU[31]) );
  OR2_X1 U46 ( .A1(n105), .A2(n745), .ZN(n668) );
  OR2_X1 U47 ( .A1(n106), .A2(n776), .ZN(n669) );
  NAND3_X1 U48 ( .A1(n107), .A2(n669), .A3(n668), .ZN(OUTALU[29]) );
  OR2_X1 U49 ( .A1(n150), .A2(n759), .ZN(n670) );
  OR2_X1 U50 ( .A1(n151), .A2(n790), .ZN(n671) );
  NAND3_X1 U51 ( .A1(n670), .A2(n671), .A3(n152), .ZN(OUTALU[15]) );
  OR2_X1 U52 ( .A1(n159), .A2(n762), .ZN(n672) );
  OR2_X1 U53 ( .A1(n160), .A2(n793), .ZN(n673) );
  NAND3_X1 U54 ( .A1(n161), .A2(n673), .A3(n672), .ZN(OUTALU[12]) );
  OR2_X1 U55 ( .A1(n123), .A2(n751), .ZN(n674) );
  OR2_X1 U56 ( .A1(n124), .A2(n782), .ZN(n675) );
  NAND3_X1 U57 ( .A1(n674), .A2(n675), .A3(n125), .ZN(OUTALU[23]) );
  OR2_X1 U58 ( .A1(n165), .A2(n764), .ZN(n676) );
  OR2_X1 U59 ( .A1(n166), .A2(n795), .ZN(n677) );
  NAND3_X1 U60 ( .A1(n676), .A2(n677), .A3(n167), .ZN(OUTALU[10]) );
  OR2_X1 U61 ( .A1(n141), .A2(n756), .ZN(n678) );
  OR2_X1 U62 ( .A1(n142), .A2(n787), .ZN(n679) );
  NAND3_X1 U63 ( .A1(n143), .A2(n679), .A3(n678), .ZN(OUTALU[18]) );
  NAND2_X1 U64 ( .A1(n104), .A2(n649), .ZN(OUTALU[2]) );
  OR2_X1 U65 ( .A1(n78), .A2(n766), .ZN(n680) );
  OR2_X1 U66 ( .A1(n79), .A2(n797), .ZN(n681) );
  NAND3_X1 U67 ( .A1(n680), .A2(n681), .A3(n80), .ZN(OUTALU[8]) );
  OR2_X1 U68 ( .A1(n108), .A2(n746), .ZN(n682) );
  OR2_X1 U69 ( .A1(n109), .A2(n777), .ZN(n683) );
  NAND3_X1 U70 ( .A1(n682), .A2(n683), .A3(n110), .ZN(OUTALU[28]) );
  NAND2_X1 U71 ( .A1(n101), .A2(n651), .ZN(OUTALU[30]) );
  BUF_X1 U72 ( .A(n74), .Z(net134765) );
  BUF_X1 U73 ( .A(n73), .Z(net134755) );
  OAI21_X1 U74 ( .B1(\Comparison[1] ), .B2(n174), .A(n175), .ZN(n74) );
  BUF_X1 U75 ( .A(n74), .Z(net134761) );
  BUF_X1 U76 ( .A(n74), .Z(net134763) );
  OR3_X1 U77 ( .A1(CODE[2]), .A2(CODE[3]), .A3(n173), .ZN(n175) );
  AND3_X1 U78 ( .A1(net131849), .A2(n684), .A3(n176), .ZN(n73) );
  BUF_X1 U79 ( .A(n73), .Z(net134759) );
  BUF_X1 U80 ( .A(n73), .Z(net134757) );
  NAND2_X1 U81 ( .A1(CODE[0]), .A2(CODE[1]), .ZN(n173) );
  NOR3_X1 U82 ( .A1(net133061), .A2(CODE[1]), .A3(n174), .ZN(n76) );
  NAND2_X1 U83 ( .A1(net131848), .A2(net133061), .ZN(\Comparison[1] ) );
  INV_X1 U84 ( .A(CODE[3]), .ZN(n684) );
  NAND2_X1 U85 ( .A1(CODE[2]), .A2(n684), .ZN(n174) );
  INV_X1 U86 ( .A(CODE[2]), .ZN(net131849) );
  NAND4_X1 U87 ( .A1(\COMPARATORout[0] ), .A2(CODE[3]), .A3(n173), .A4(
        net131849), .ZN(n172) );
  NOR2_X1 U88 ( .A1(n174), .A2(n173), .ZN(n75) );
  INV_X1 U89 ( .A(CODE[1]), .ZN(net131848) );
  INV_X1 U90 ( .A(DATA2[4]), .ZN(net131855) );
  AOI21_X1 U91 ( .B1(net134775), .B2(net131855), .A(net134793), .ZN(n90) );
  AOI221_X1 U92 ( .B1(net134767), .B2(net131887), .C1(DATA1[4]), .C2(net134783), .A(net134785), .ZN(n91) );
  BUF_X1 U93 ( .A(n77), .Z(net134785) );
  BUF_X1 U94 ( .A(n76), .Z(net134783) );
  INV_X1 U95 ( .A(DATA1[4]), .ZN(net131887) );
  BUF_X1 U96 ( .A(n75), .Z(net134767) );
  BUF_X1 U97 ( .A(n77), .Z(net134793) );
  BUF_X1 U98 ( .A(n75), .Z(net134775) );
  INV_X1 U99 ( .A(n804), .ZN(n685) );
  CLKBUF_X1 U100 ( .A(DATA2[27]), .Z(n686) );
  CLKBUF_X1 U101 ( .A(DATA2[8]), .Z(n687) );
  CLKBUF_X1 U102 ( .A(DATA2[20]), .Z(n688) );
  CLKBUF_X1 U103 ( .A(DATA2[11]), .Z(n689) );
  CLKBUF_X1 U104 ( .A(DATA2[19]), .Z(n691) );
  CLKBUF_X1 U105 ( .A(DATA2[9]), .Z(n692) );
  CLKBUF_X1 U106 ( .A(DATA2[14]), .Z(n693) );
  CLKBUF_X1 U107 ( .A(DATA2[21]), .Z(n694) );
  CLKBUF_X1 U108 ( .A(DATA2[30]), .Z(n695) );
  NAND2_X1 U109 ( .A1(n137), .A2(n650), .ZN(OUTALU[1]) );
  CLKBUF_X1 U110 ( .A(DATA2[6]), .Z(n696) );
  CLKBUF_X1 U111 ( .A(DATA2[26]), .Z(n697) );
  CLKBUF_X1 U112 ( .A(DATA2[29]), .Z(n698) );
  CLKBUF_X1 U113 ( .A(DATA2[12]), .Z(n700) );
  CLKBUF_X1 U114 ( .A(DATA2[28]), .Z(n701) );
  CLKBUF_X1 U115 ( .A(DATA2[24]), .Z(n702) );
  CLKBUF_X1 U116 ( .A(DATA2[25]), .Z(n703) );
  CLKBUF_X1 U117 ( .A(DATA2[23]), .Z(n705) );
  CLKBUF_X1 U118 ( .A(DATA2[10]), .Z(n706) );
  CLKBUF_X1 U119 ( .A(DATA2[16]), .Z(n707) );
  CLKBUF_X1 U120 ( .A(DATA2[18]), .Z(n708) );
  OR2_X1 U121 ( .A1(n156), .A2(n761), .ZN(n709) );
  OR2_X1 U122 ( .A1(n157), .A2(n792), .ZN(n710) );
  NAND3_X1 U123 ( .A1(n158), .A2(n710), .A3(n709), .ZN(OUTALU[13]) );
  CLKBUF_X1 U124 ( .A(DATA2[17]), .Z(n711) );
  NAND3_X1 U125 ( .A1(n733), .A2(n734), .A3(n735), .ZN(OUTALU[0]) );
  OR2_X1 U126 ( .A1(n99), .A2(n744), .ZN(n713) );
  OR2_X1 U127 ( .A1(n100), .A2(n775), .ZN(n714) );
  OR2_X1 U128 ( .A1(n70), .A2(n765), .ZN(n715) );
  OR2_X1 U129 ( .A1(n71), .A2(n796), .ZN(n716) );
  NAND3_X1 U130 ( .A1(n72), .A2(n716), .A3(n715), .ZN(OUTALU[9]) );
  OR2_X1 U131 ( .A1(n144), .A2(n757), .ZN(n717) );
  OR2_X1 U132 ( .A1(n145), .A2(n788), .ZN(n718) );
  NAND3_X1 U133 ( .A1(n717), .A2(n718), .A3(n146), .ZN(OUTALU[17]) );
  OR2_X1 U134 ( .A1(n93), .A2(n770), .ZN(n719) );
  OR2_X1 U135 ( .A1(n94), .A2(n801), .ZN(n720) );
  NAND3_X1 U136 ( .A1(n95), .A2(n720), .A3(n719), .ZN(OUTALU[3]) );
  OR2_X1 U137 ( .A1(n117), .A2(n749), .ZN(n721) );
  OR2_X1 U138 ( .A1(n118), .A2(n780), .ZN(n722) );
  NAND3_X1 U139 ( .A1(n119), .A2(n722), .A3(n721), .ZN(OUTALU[25]) );
  OR2_X1 U140 ( .A1(n162), .A2(n763), .ZN(n723) );
  OR2_X1 U141 ( .A1(n163), .A2(n794), .ZN(n724) );
  NAND3_X1 U142 ( .A1(n164), .A2(n724), .A3(n723), .ZN(OUTALU[11]) );
  OR2_X1 U143 ( .A1(n126), .A2(n752), .ZN(n725) );
  OR2_X1 U144 ( .A1(n127), .A2(n783), .ZN(n726) );
  OR2_X1 U145 ( .A1(n102), .A2(n771), .ZN(n727) );
  OR2_X1 U146 ( .A1(n103), .A2(n802), .ZN(n728) );
  OR2_X1 U147 ( .A1(n135), .A2(n772), .ZN(n729) );
  OR2_X1 U148 ( .A1(n136), .A2(n803), .ZN(n730) );
  OR2_X1 U149 ( .A1(n84), .A2(n768), .ZN(n731) );
  OR2_X1 U150 ( .A1(n85), .A2(n799), .ZN(n732) );
  NAND3_X1 U151 ( .A1(n86), .A2(n732), .A3(n731), .ZN(OUTALU[6]) );
  NAND2_X1 U152 ( .A1(SHIFTERout[0]), .A2(net134759), .ZN(n733) );
  NAND2_X1 U153 ( .A1(ADDERout[0]), .A2(net134761), .ZN(n734) );
  INV_X1 U154 ( .A(n169), .ZN(n735) );
  BUF_X1 U155 ( .A(n75), .Z(net134771) );
  BUF_X1 U156 ( .A(n75), .Z(net134769) );
  BUF_X1 U157 ( .A(n75), .Z(net134773) );
  BUF_X1 U158 ( .A(n77), .Z(net134789) );
  BUF_X1 U159 ( .A(n77), .Z(net134791) );
  BUF_X1 U160 ( .A(n77), .Z(net134787) );
  AOI22_X1 U161 ( .A1(SHIFTERout[14]), .A2(net134759), .B1(ADDERout[14]), .B2(
        net134761), .ZN(n155) );
  AOI22_X1 U162 ( .A1(SHIFTERout[15]), .A2(net134759), .B1(ADDERout[15]), .B2(
        net134761), .ZN(n152) );
  AOI22_X1 U163 ( .A1(SHIFTERout[10]), .A2(net134759), .B1(ADDERout[10]), .B2(
        net134761), .ZN(n167) );
  AOI22_X1 U164 ( .A1(SHIFTERout[19]), .A2(net134757), .B1(ADDERout[19]), .B2(
        net134761), .ZN(n140) );
  AOI221_X1 U165 ( .B1(net134769), .B2(n755), .C1(DATA1[19]), .C2(net134779), 
        .A(net134787), .ZN(n139) );
  AOI221_X1 U166 ( .B1(net134767), .B2(n746), .C1(DATA1[28]), .C2(net134781), 
        .A(net134785), .ZN(n109) );
  AOI221_X1 U167 ( .B1(net134769), .B2(n765), .C1(net134783), .C2(DATA1[9]), 
        .A(net134787), .ZN(n71) );
  AOI221_X1 U168 ( .B1(net134769), .B2(n772), .C1(DATA1[1]), .C2(net134779), 
        .A(net134787), .ZN(n136) );
  AOI221_X1 U169 ( .B1(net134771), .B2(n761), .C1(DATA1[13]), .C2(net134779), 
        .A(net134789), .ZN(n157) );
  AOI221_X1 U170 ( .B1(net134767), .B2(n770), .C1(DATA1[3]), .C2(net134783), 
        .A(net134785), .ZN(n94) );
  AOI221_X1 U171 ( .B1(net134769), .B2(n749), .C1(DATA1[25]), .C2(net134781), 
        .A(net134787), .ZN(n118) );
  AOI221_X1 U172 ( .B1(net134769), .B2(n751), .C1(DATA1[23]), .C2(net134781), 
        .A(net134787), .ZN(n124) );
  AOI221_X1 U173 ( .B1(net134767), .B2(n768), .C1(DATA1[6]), .C2(net134783), 
        .A(net134785), .ZN(n85) );
  AOI221_X1 U174 ( .B1(net134767), .B2(n766), .C1(DATA1[8]), .C2(net134783), 
        .A(net134785), .ZN(n79) );
  AOI221_X1 U175 ( .B1(net134771), .B2(n763), .C1(DATA1[11]), .C2(net134779), 
        .A(net134789), .ZN(n163) );
  AOI221_X1 U176 ( .B1(net134771), .B2(n760), .C1(DATA1[14]), .C2(net134779), 
        .A(net134789), .ZN(n154) );
  AOI221_X1 U177 ( .B1(net134771), .B2(n759), .C1(DATA1[15]), .C2(net134779), 
        .A(net134789), .ZN(n151) );
  AOI221_X1 U178 ( .B1(net134771), .B2(n757), .C1(DATA1[17]), .C2(net134779), 
        .A(net134789), .ZN(n145) );
  AOI221_X1 U179 ( .B1(net134769), .B2(n756), .C1(DATA1[18]), .C2(net134779), 
        .A(net134787), .ZN(n142) );
  AOI221_X1 U180 ( .B1(net134769), .B2(n752), .C1(DATA1[22]), .C2(net134781), 
        .A(net134787), .ZN(n127) );
  AOI221_X1 U181 ( .B1(net134767), .B2(n745), .C1(DATA1[29]), .C2(net134781), 
        .A(net134785), .ZN(n106) );
  AOI221_X1 U182 ( .B1(net134767), .B2(n743), .C1(DATA1[31]), .C2(net134783), 
        .A(net134785), .ZN(n97) );
  BUF_X1 U183 ( .A(n76), .Z(net134779) );
  BUF_X1 U184 ( .A(n76), .Z(net134781) );
  INV_X1 U185 ( .A(DATA1[30]), .ZN(n744) );
  INV_X1 U186 ( .A(DATA1[29]), .ZN(n745) );
  INV_X1 U187 ( .A(DATA1[25]), .ZN(n749) );
  INV_X1 U188 ( .A(DATA1[1]), .ZN(n772) );
  INV_X1 U189 ( .A(DATA1[22]), .ZN(n752) );
  INV_X1 U190 ( .A(DATA1[26]), .ZN(n748) );
  INV_X1 U191 ( .A(DATA1[23]), .ZN(n751) );
  INV_X1 U192 ( .A(DATA1[31]), .ZN(n743) );
  INV_X1 U193 ( .A(DATA1[28]), .ZN(n746) );
  INV_X1 U194 ( .A(DATA1[13]), .ZN(n761) );
  INV_X1 U195 ( .A(DATA1[8]), .ZN(n766) );
  INV_X1 U196 ( .A(DATA1[19]), .ZN(n755) );
  INV_X1 U197 ( .A(DATA1[6]), .ZN(n768) );
  INV_X1 U198 ( .A(DATA1[15]), .ZN(n759) );
  INV_X1 U199 ( .A(DATA1[17]), .ZN(n757) );
  INV_X1 U200 ( .A(DATA1[18]), .ZN(n756) );
  INV_X1 U201 ( .A(DATA1[21]), .ZN(n753) );
  INV_X1 U202 ( .A(DATA1[24]), .ZN(n750) );
  INV_X1 U203 ( .A(DATA1[12]), .ZN(n762) );
  INV_X1 U204 ( .A(DATA1[7]), .ZN(n767) );
  INV_X1 U205 ( .A(DATA1[14]), .ZN(n760) );
  INV_X1 U206 ( .A(DATA1[27]), .ZN(n747) );
  INV_X1 U207 ( .A(DATA1[9]), .ZN(n765) );
  INV_X1 U208 ( .A(DATA1[11]), .ZN(n763) );
  INV_X1 U210 ( .A(DATA1[3]), .ZN(n770) );
  INV_X1 U211 ( .A(DATA1[0]), .ZN(n773) );
  INV_X1 U212 ( .A(n711), .ZN(n788) );
  INV_X1 U213 ( .A(n687), .ZN(n797) );
  INV_X1 U214 ( .A(n686), .ZN(n778) );
  INV_X1 U215 ( .A(n697), .ZN(n779) );
  INV_X1 U216 ( .A(DATA2[1]), .ZN(n803) );
  INV_X1 U217 ( .A(n663), .ZN(n802) );
  INV_X1 U218 ( .A(DATA2[3]), .ZN(n801) );
  AOI221_X1 U219 ( .B1(net134769), .B2(n758), .C1(DATA1[16]), .C2(net134779), 
        .A(net134787), .ZN(n148) );
  AOI221_X1 U220 ( .B1(net134769), .B2(n754), .C1(DATA1[20]), .C2(net134781), 
        .A(net134787), .ZN(n133) );
  AOI221_X1 U221 ( .B1(net134767), .B2(n769), .C1(DATA1[5]), .C2(net134783), 
        .A(net134785), .ZN(n88) );
  AOI221_X1 U222 ( .B1(net134767), .B2(n771), .C1(DATA1[2]), .C2(net134781), 
        .A(net134785), .ZN(n103) );
  AOI221_X1 U223 ( .B1(net134771), .B2(n764), .C1(DATA1[10]), .C2(net134779), 
        .A(net134789), .ZN(n166) );
  AOI21_X1 U224 ( .B1(net134777), .B2(n804), .A(net134795), .ZN(n170) );
  AOI221_X1 U225 ( .B1(net134771), .B2(n773), .C1(DATA1[0]), .C2(net134779), 
        .A(net134789), .ZN(n171) );
  AOI21_X1 U226 ( .B1(net134773), .B2(n778), .A(net134791), .ZN(n111) );
  AOI21_X1 U227 ( .B1(net134773), .B2(n791), .A(net134791), .ZN(n153) );
  AOI21_X1 U228 ( .B1(net134771), .B2(n783), .A(net134789), .ZN(n126) );
  AOI21_X1 U229 ( .B1(net134771), .B2(n786), .A(net134789), .ZN(n138) );
  AOI21_X1 U230 ( .B1(net134773), .B2(n782), .A(net134791), .ZN(n123) );
  AOI21_X1 U231 ( .B1(net134773), .B2(n787), .A(net134791), .ZN(n141) );
  AOI21_X1 U232 ( .B1(net134773), .B2(n780), .A(net134791), .ZN(n117) );
  AOI21_X1 U233 ( .B1(net134773), .B2(n777), .A(net134791), .ZN(n108) );
  AOI21_X1 U234 ( .B1(net134775), .B2(n792), .A(net134793), .ZN(n156) );
  AOI21_X1 U235 ( .B1(net134773), .B2(n788), .A(net134791), .ZN(n144) );
  AOI21_X1 U236 ( .B1(net134773), .B2(n779), .A(net134791), .ZN(n114) );
  AOI21_X1 U237 ( .B1(net134775), .B2(n776), .A(net134793), .ZN(n105) );
  AOI21_X1 U238 ( .B1(net134775), .B2(n775), .A(net134793), .ZN(n99) );
  AOI21_X1 U239 ( .B1(net134771), .B2(n784), .A(net134789), .ZN(n129) );
  AOI21_X1 U240 ( .B1(net134775), .B2(n794), .A(net134793), .ZN(n162) );
  AOI21_X1 U241 ( .B1(net134777), .B2(n796), .A(net134795), .ZN(n70) );
  AOI21_X1 U242 ( .B1(net134775), .B2(n799), .A(net134793), .ZN(n84) );
  AOI21_X1 U243 ( .B1(net134773), .B2(n781), .A(net134791), .ZN(n120) );
  AOI21_X1 U244 ( .B1(net134777), .B2(n797), .A(net134793), .ZN(n78) );
  AOI21_X1 U245 ( .B1(net134775), .B2(n793), .A(net134793), .ZN(n159) );
  AOI21_X1 U246 ( .B1(net134775), .B2(n801), .A(net134793), .ZN(n93) );
  AOI21_X1 U247 ( .B1(net134775), .B2(n798), .A(net134793), .ZN(n81) );
  AOI21_X1 U248 ( .B1(net134775), .B2(n774), .A(net134793), .ZN(n96) );
  AOI21_X1 U249 ( .B1(net134773), .B2(n802), .A(net134791), .ZN(n102) );
  AOI21_X1 U250 ( .B1(net134771), .B2(n803), .A(net134789), .ZN(n135) );
  AOI21_X1 U251 ( .B1(net134775), .B2(n790), .A(net134791), .ZN(n150) );
  AOI21_X1 U252 ( .B1(net134777), .B2(n795), .A(net134793), .ZN(n165) );
  INV_X1 U253 ( .A(DATA1[2]), .ZN(n771) );
  INV_X1 U254 ( .A(DATA1[10]), .ZN(n764) );
  INV_X1 U255 ( .A(n693), .ZN(n791) );
  INV_X1 U256 ( .A(n704), .ZN(n792) );
  INV_X1 U257 ( .A(n700), .ZN(n793) );
  AOI22_X1 U258 ( .A1(SHIFTERout[26]), .A2(net134757), .B1(ADDERout[26]), .B2(
        net134763), .ZN(n116) );
  INV_X1 U259 ( .A(n695), .ZN(n775) );
  AOI22_X1 U260 ( .A1(SHIFTERout[18]), .A2(net134757), .B1(ADDERout[18]), .B2(
        net134761), .ZN(n143) );
  OAI221_X1 U261 ( .B1(n170), .B2(n773), .C1(n171), .C2(n804), .A(n172), .ZN(
        n169) );
  AOI22_X1 U262 ( .A1(SHIFTERout[24]), .A2(net134757), .B1(ADDERout[24]), .B2(
        net134763), .ZN(n122) );
  AOI22_X1 U263 ( .A1(SHIFTERout[31]), .A2(net134755), .B1(ADDERout[31]), .B2(
        net134765), .ZN(n98) );
  CLKBUF_X1 U264 ( .A(DATA2[22]), .Z(n736) );
  OR2_X1 U265 ( .A1(n147), .A2(n758), .ZN(n737) );
  OR2_X1 U266 ( .A1(n148), .A2(n789), .ZN(n738) );
  NAND3_X1 U267 ( .A1(n149), .A2(n738), .A3(n737), .ZN(OUTALU[16]) );
  AOI21_X1 U268 ( .B1(net134773), .B2(n789), .A(net134791), .ZN(n147) );
  INV_X1 U269 ( .A(DATA1[16]), .ZN(n758) );
  AOI22_X1 U270 ( .A1(SHIFTERout[11]), .A2(net134759), .B1(ADDERout[11]), .B2(
        net134761), .ZN(n164) );
  OR2_X1 U271 ( .A1(n132), .A2(n754), .ZN(n739) );
  OR2_X1 U272 ( .A1(n133), .A2(n785), .ZN(n740) );
  NAND3_X1 U273 ( .A1(n739), .A2(n740), .A3(n134), .ZN(OUTALU[20]) );
  AOI21_X1 U274 ( .B1(net134773), .B2(n785), .A(net134791), .ZN(n132) );
  INV_X1 U275 ( .A(DATA1[20]), .ZN(n754) );
  AOI22_X1 U276 ( .A1(SHIFTERout[25]), .A2(net134757), .B1(ADDERout[25]), .B2(
        net134763), .ZN(n119) );
  AOI22_X1 U277 ( .A1(SHIFTERout[22]), .A2(net134757), .B1(ADDERout[22]), .B2(
        net134763), .ZN(n128) );
  AOI22_X1 U278 ( .A1(SHIFTERout[23]), .A2(net134757), .B1(ADDERout[23]), .B2(
        net134763), .ZN(n125) );
  AOI22_X1 U279 ( .A1(SHIFTERout[9]), .A2(net134755), .B1(ADDERout[9]), .B2(
        net134765), .ZN(n72) );
  INV_X1 U280 ( .A(n698), .ZN(n776) );
  INV_X1 U281 ( .A(n708), .ZN(n787) );
  OAI221_X1 U282 ( .B1(n138), .B2(n755), .C1(n139), .C2(n786), .A(n140), .ZN(
        OUTALU[19]) );
  AOI22_X1 U283 ( .A1(SHIFTERout[17]), .A2(net134757), .B1(ADDERout[17]), .B2(
        net134761), .ZN(n146) );
  OR2_X1 U284 ( .A1(n87), .A2(n769), .ZN(n741) );
  OR2_X1 U285 ( .A1(n88), .A2(n800), .ZN(n742) );
  AOI21_X1 U286 ( .B1(net134775), .B2(n800), .A(net134793), .ZN(n87) );
  INV_X1 U287 ( .A(DATA1[5]), .ZN(n769) );
  INV_X1 U288 ( .A(DATA2[5]), .ZN(n800) );
  INV_X1 U289 ( .A(n692), .ZN(n796) );
  AOI22_X1 U290 ( .A1(SHIFTERout[16]), .A2(net134759), .B1(ADDERout[16]), .B2(
        net134761), .ZN(n149) );
  INV_X1 U291 ( .A(n691), .ZN(n786) );
  AOI22_X1 U292 ( .A1(SHIFTERout[20]), .A2(net134757), .B1(ADDERout[20]), .B2(
        net134763), .ZN(n134) );
  INV_X1 U293 ( .A(DATA2[31]), .ZN(n774) );
  OAI221_X1 U294 ( .B1(n153), .B2(n760), .C1(n154), .C2(n791), .A(n155), .ZN(
        OUTALU[14]) );
  INV_X1 U295 ( .A(n690), .ZN(n798) );
  AOI22_X1 U296 ( .A1(SHIFTERout[6]), .A2(net134755), .B1(ADDERout[6]), .B2(
        net134765), .ZN(n86) );
  AOI22_X1 U297 ( .A1(SHIFTERout[30]), .A2(net134755), .B1(ADDERout[30]), .B2(
        net134763), .ZN(n101) );
  INV_X1 U298 ( .A(n694), .ZN(n784) );
  AOI22_X1 U299 ( .A1(SHIFTERout[13]), .A2(net134759), .B1(ADDERout[13]), .B2(
        net134761), .ZN(n158) );
  AOI22_X1 U300 ( .A1(SHIFTERout[12]), .A2(net134759), .B1(ADDERout[12]), .B2(
        net134761), .ZN(n161) );
  AOI22_X1 U301 ( .A1(SHIFTERout[2]), .A2(net134755), .B1(ADDERout[2]), .B2(
        net134763), .ZN(n104) );
  INV_X1 U302 ( .A(n699), .ZN(n790) );
  OAI221_X1 U303 ( .B1(n81), .B2(n767), .C1(n82), .C2(n798), .A(n83), .ZN(
        OUTALU[7]) );
  AOI22_X1 U304 ( .A1(SHIFTERout[7]), .A2(net134755), .B1(ADDERout[7]), .B2(
        net134765), .ZN(n83) );
  INV_X1 U305 ( .A(DATA2[0]), .ZN(n804) );
  AOI22_X1 U306 ( .A1(SHIFTERout[29]), .A2(net134755), .B1(ADDERout[29]), .B2(
        net134763), .ZN(n107) );
  INV_X1 U307 ( .A(n707), .ZN(n789) );
  INV_X1 U308 ( .A(n688), .ZN(n785) );
  INV_X1 U309 ( .A(n703), .ZN(n780) );
  OAI221_X1 U310 ( .B1(n114), .B2(n748), .C1(n115), .C2(n779), .A(n116), .ZN(
        OUTALU[26]) );
  INV_X1 U311 ( .A(n689), .ZN(n794) );
  INV_X1 U312 ( .A(n705), .ZN(n782) );
  INV_X1 U313 ( .A(n702), .ZN(n781) );
  AOI22_X1 U314 ( .A1(SHIFTERout[27]), .A2(net134757), .B1(ADDERout[27]), .B2(
        net134763), .ZN(n113) );
  OAI221_X1 U315 ( .B1(n111), .B2(n747), .C1(n112), .C2(n778), .A(n113), .ZN(
        OUTALU[27]) );
  INV_X1 U316 ( .A(n706), .ZN(n795) );
  INV_X1 U317 ( .A(n696), .ZN(n799) );
  INV_X1 U318 ( .A(n701), .ZN(n777) );
  AOI22_X1 U319 ( .A1(SHIFTERout[28]), .A2(net134755), .B1(ADDERout[28]), .B2(
        net134763), .ZN(n110) );
  INV_X1 U320 ( .A(n736), .ZN(n783) );
  CLKBUF_X1 U321 ( .A(n77), .Z(net134795) );
  CLKBUF_X1 U322 ( .A(n75), .Z(net134777) );
endmodule


module reg_6 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n93, n94, n95, n96, n97, n98, n99, n102, net134801, net134799,
         net134797, net134807, net134805, net134803, n35, n34, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204;

  DFF_X1 \temp_reg[27]  ( .D(n71), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n72), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[24]  ( .D(n74), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[22]  ( .D(n76), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n77), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[18]  ( .D(n80), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n81), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n82), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n83), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n84), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[11]  ( .D(n87), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n88), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[8]  ( .D(n90), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n91), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n102), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n93), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n94), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[2]  ( .D(n96), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[0]  ( .D(n98), .CK(clock), .Q(o[0]), .QN(n36) );
  DFF_X1 \temp_reg[23]  ( .D(n75), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[25]  ( .D(n73), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[3]  ( .D(n95), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[13]  ( .D(n85), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[1]  ( .D(n97), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[9]  ( .D(n89), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[20]  ( .D(n78), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n79), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[12]  ( .D(n86), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[28]  ( .D(n70), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[31]  ( .D(n99), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[29]  ( .D(n69), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[30]  ( .D(n68), .CK(clock), .Q(o[30]), .QN(n66) );
  BUF_X1 U3 ( .A(n35), .Z(net134807) );
  BUF_X1 U4 ( .A(n34), .Z(net134801) );
  BUF_X1 U5 ( .A(n35), .Z(net134805) );
  BUF_X1 U6 ( .A(n34), .Z(net134799) );
  BUF_X1 U7 ( .A(n35), .Z(net134803) );
  BUF_X1 U8 ( .A(n34), .Z(net134797) );
  OAI22_X1 U9 ( .A1(n176), .A2(n34), .B1(n35), .B2(n45), .ZN(n89) );
  OAI22_X1 U10 ( .A1(n202), .A2(n34), .B1(n35), .B2(n42), .ZN(n102) );
  OAI22_X1 U11 ( .A1(n180), .A2(n34), .B1(n35), .B2(n49), .ZN(n85) );
  OAI22_X1 U12 ( .A1(n185), .A2(n34), .B1(n35), .B2(n52), .ZN(n82) );
  OAI22_X1 U13 ( .A1(n190), .A2(n34), .B1(n35), .B2(n63), .ZN(n71) );
  OAI22_X1 U14 ( .A1(n191), .A2(n34), .B1(n35), .B2(n62), .ZN(n72) );
  OAI22_X1 U15 ( .A1(n184), .A2(n34), .B1(n35), .B2(n53), .ZN(n81) );
  OAI22_X1 U16 ( .A1(n188), .A2(n34), .B1(n35), .B2(n57), .ZN(n77) );
  OAI22_X1 U17 ( .A1(n172), .A2(n34), .B1(n35), .B2(n40), .ZN(n94) );
  INV_X1 U18 ( .A(i[4]), .ZN(n172) );
  OR2_X1 U19 ( .A1(reset), .A2(load), .ZN(n35) );
  NAND2_X1 U20 ( .A1(load), .A2(n173), .ZN(n34) );
  INV_X1 U21 ( .A(reset), .ZN(n173) );
  OAI22_X1 U22 ( .A1(net134799), .A2(n178), .B1(net134805), .B2(n51), .ZN(n83)
         );
  INV_X1 U23 ( .A(i[10]), .ZN(n175) );
  OAI22_X1 U24 ( .A1(net134801), .A2(n194), .B1(net134807), .B2(n67), .ZN(n99)
         );
  OAI22_X1 U25 ( .A1(net134797), .A2(n193), .B1(net134803), .B2(n60), .ZN(n74)
         );
  INV_X1 U26 ( .A(i[28]), .ZN(n197) );
  INV_X1 U27 ( .A(i[27]), .ZN(n190) );
  OAI22_X1 U28 ( .A1(net134801), .A2(n199), .B1(net134807), .B2(n43), .ZN(n91)
         );
  INV_X1 U29 ( .A(i[7]), .ZN(n199) );
  OAI22_X1 U30 ( .A1(net134799), .A2(n179), .B1(net134805), .B2(n50), .ZN(n84)
         );
  OAI22_X1 U31 ( .A1(net134799), .A2(n181), .B1(net134805), .B2(n48), .ZN(n86)
         );
  OAI22_X1 U32 ( .A1(n198), .A2(net134801), .B1(net134807), .B2(n36), .ZN(n98)
         );
  INV_X1 U33 ( .A(i[0]), .ZN(n198) );
  OAI22_X1 U34 ( .A1(net134799), .A2(n183), .B1(net134805), .B2(n54), .ZN(n80)
         );
  OAI22_X1 U35 ( .A1(n192), .A2(net134797), .B1(net134803), .B2(n61), .ZN(n73)
         );
  INV_X1 U36 ( .A(i[17]), .ZN(n184) );
  INV_X1 U37 ( .A(i[12]), .ZN(n181) );
  OAI22_X1 U38 ( .A1(net134797), .A2(n197), .B1(net134803), .B2(n64), .ZN(n70)
         );
  OAI22_X1 U39 ( .A1(net134797), .A2(n195), .B1(net134803), .B2(n66), .ZN(n68)
         );
  INV_X1 U40 ( .A(i[16]), .ZN(n185) );
  INV_X1 U41 ( .A(i[13]), .ZN(n180) );
  INV_X1 U42 ( .A(i[5]), .ZN(n204) );
  INV_X1 U43 ( .A(i[24]), .ZN(n193) );
  INV_X1 U44 ( .A(i[14]), .ZN(n179) );
  INV_X1 U45 ( .A(i[9]), .ZN(n176) );
  OAI22_X1 U46 ( .A1(n203), .A2(net134801), .B1(net134807), .B2(n37), .ZN(n97)
         );
  INV_X1 U47 ( .A(i[31]), .ZN(n194) );
  OAI22_X1 U48 ( .A1(net134797), .A2(n196), .B1(net134803), .B2(n65), .ZN(n69)
         );
  INV_X1 U49 ( .A(i[15]), .ZN(n178) );
  OAI22_X1 U50 ( .A1(net134799), .A2(n177), .B1(net134805), .B2(n44), .ZN(n90)
         );
  OAI22_X1 U51 ( .A1(net134797), .A2(n187), .B1(net134803), .B2(n58), .ZN(n76)
         );
  OAI22_X1 U52 ( .A1(n200), .A2(net134801), .B1(net134807), .B2(n39), .ZN(n95)
         );
  OAI22_X1 U53 ( .A1(net134799), .A2(n175), .B1(net134805), .B2(n46), .ZN(n88)
         );
  INV_X1 U54 ( .A(i[18]), .ZN(n183) );
  INV_X1 U55 ( .A(i[21]), .ZN(n188) );
  OAI22_X1 U56 ( .A1(net134797), .A2(n186), .B1(net134803), .B2(n59), .ZN(n75)
         );
  INV_X1 U57 ( .A(i[23]), .ZN(n186) );
  OAI22_X1 U58 ( .A1(n204), .A2(net134801), .B1(net134807), .B2(n41), .ZN(n93)
         );
  INV_X1 U59 ( .A(i[3]), .ZN(n200) );
  INV_X1 U60 ( .A(i[30]), .ZN(n195) );
  INV_X1 U61 ( .A(i[26]), .ZN(n191) );
  OAI22_X1 U62 ( .A1(n174), .A2(net134799), .B1(net134805), .B2(n47), .ZN(n87)
         );
  INV_X1 U63 ( .A(i[11]), .ZN(n174) );
  INV_X1 U64 ( .A(i[22]), .ZN(n187) );
  INV_X1 U65 ( .A(i[25]), .ZN(n192) );
  OAI22_X1 U66 ( .A1(n189), .A2(net134797), .B1(net134803), .B2(n56), .ZN(n78)
         );
  INV_X1 U67 ( .A(i[20]), .ZN(n189) );
  INV_X1 U68 ( .A(i[8]), .ZN(n177) );
  INV_X1 U69 ( .A(i[6]), .ZN(n202) );
  OAI22_X1 U70 ( .A1(n201), .A2(net134801), .B1(net134807), .B2(n38), .ZN(n96)
         );
  INV_X1 U71 ( .A(i[2]), .ZN(n201) );
  OAI22_X1 U72 ( .A1(net134799), .A2(n182), .B1(net134805), .B2(n55), .ZN(n79)
         );
  INV_X1 U73 ( .A(i[19]), .ZN(n182) );
  INV_X1 U74 ( .A(i[1]), .ZN(n203) );
  INV_X1 U75 ( .A(i[29]), .ZN(n196) );
endmodule


module reg_5 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n215), .Z(n177) );
  BUF_X1 U4 ( .A(n215), .Z(n176) );
  BUF_X1 U5 ( .A(n215), .Z(n178) );
  BUF_X1 U6 ( .A(n216), .Z(n179) );
  BUF_X1 U7 ( .A(n216), .Z(n180) );
  BUF_X1 U8 ( .A(n216), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n215) );
  OAI22_X1 U10 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U12 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n213) );
  OAI22_X1 U14 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U16 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U18 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U20 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U22 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U24 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U26 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U28 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n205) );
  OAI22_X1 U30 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U32 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U34 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U36 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U38 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U40 ( .A1(n180), .A2(n51), .B1(n177), .B2(n199), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n199) );
  OAI22_X1 U42 ( .A1(n180), .A2(n52), .B1(n177), .B2(n198), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n198) );
  OAI22_X1 U44 ( .A1(n180), .A2(n53), .B1(n177), .B2(n197), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n197) );
  OAI22_X1 U46 ( .A1(n180), .A2(n54), .B1(n177), .B2(n196), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n196) );
  OAI22_X1 U48 ( .A1(n180), .A2(n55), .B1(n177), .B2(n195), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n195) );
  OAI22_X1 U50 ( .A1(n179), .A2(n56), .B1(n176), .B2(n194), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n194) );
  OAI22_X1 U52 ( .A1(n179), .A2(n57), .B1(n176), .B2(n193), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n193) );
  OAI22_X1 U54 ( .A1(n179), .A2(n58), .B1(n176), .B2(n192), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n192) );
  OAI22_X1 U56 ( .A1(n179), .A2(n59), .B1(n176), .B2(n191), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n191) );
  OAI22_X1 U58 ( .A1(n179), .A2(n60), .B1(n176), .B2(n190), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n190) );
  OAI22_X1 U60 ( .A1(n179), .A2(n61), .B1(n176), .B2(n189), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n189) );
  OAI22_X1 U62 ( .A1(n179), .A2(n62), .B1(n176), .B2(n188), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n188) );
  OAI22_X1 U64 ( .A1(n179), .A2(n63), .B1(n176), .B2(n187), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n187) );
  OAI22_X1 U66 ( .A1(n179), .A2(n64), .B1(n176), .B2(n186), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n186) );
  OAI22_X1 U68 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U70 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U72 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n183) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n216) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module reg_4 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n215), .Z(n177) );
  BUF_X1 U4 ( .A(n215), .Z(n176) );
  BUF_X1 U5 ( .A(n215), .Z(n178) );
  BUF_X1 U6 ( .A(n216), .Z(n179) );
  BUF_X1 U7 ( .A(n216), .Z(n180) );
  BUF_X1 U8 ( .A(n216), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n215) );
  OAI22_X1 U10 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U12 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n213) );
  OAI22_X1 U14 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U16 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U18 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U20 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U22 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U24 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U26 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U28 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n205) );
  OAI22_X1 U30 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U32 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U34 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U36 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U38 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U40 ( .A1(n180), .A2(n51), .B1(n177), .B2(n199), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n199) );
  OAI22_X1 U42 ( .A1(n180), .A2(n52), .B1(n177), .B2(n198), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n198) );
  OAI22_X1 U44 ( .A1(n180), .A2(n53), .B1(n177), .B2(n197), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n197) );
  OAI22_X1 U46 ( .A1(n180), .A2(n54), .B1(n177), .B2(n196), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n196) );
  OAI22_X1 U48 ( .A1(n180), .A2(n55), .B1(n177), .B2(n195), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n195) );
  OAI22_X1 U50 ( .A1(n179), .A2(n56), .B1(n176), .B2(n194), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n194) );
  OAI22_X1 U52 ( .A1(n179), .A2(n57), .B1(n176), .B2(n193), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n193) );
  OAI22_X1 U54 ( .A1(n179), .A2(n58), .B1(n176), .B2(n192), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n192) );
  OAI22_X1 U56 ( .A1(n179), .A2(n59), .B1(n176), .B2(n191), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n191) );
  OAI22_X1 U58 ( .A1(n179), .A2(n60), .B1(n176), .B2(n190), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n190) );
  OAI22_X1 U60 ( .A1(n179), .A2(n61), .B1(n176), .B2(n189), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n189) );
  OAI22_X1 U62 ( .A1(n179), .A2(n62), .B1(n176), .B2(n188), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n188) );
  OAI22_X1 U64 ( .A1(n179), .A2(n63), .B1(n176), .B2(n187), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n187) );
  OAI22_X1 U66 ( .A1(n179), .A2(n64), .B1(n176), .B2(n186), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n186) );
  OAI22_X1 U68 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U70 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U72 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n183) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n216) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module executeUnit_M32_C4 ( clock, reset, en3, Mux1Sel, Mux2Sel, ALUCODE, 
        OUT1RF, OUT2RF, IMMEDIATE, NPCFromDecode, AddressWfromDecode, 
        ALUtoMEMORY, OUT2RFtoMEMORY, AddressWtoMEMORY );
  input [3:0] ALUCODE;
  input [31:0] OUT1RF;
  input [31:0] OUT2RF;
  input [31:0] IMMEDIATE;
  input [31:0] NPCFromDecode;
  input [31:0] AddressWfromDecode;
  output [31:0] ALUtoMEMORY;
  output [31:0] OUT2RFtoMEMORY;
  output [31:0] AddressWtoMEMORY;
  input clock, reset, en3, Mux1Sel, Mux2Sel;

  wire   [31:0] MUX2out;
  wire   [31:0] MUXNPCout;
  wire   [31:0] MUXWITH4out;
  wire   [31:0] ALUout;

  Mux21_4 MUX ( .a(OUT2RF), .b(IMMEDIATE), .sel(Mux2Sel), .y(MUX2out) );
  Mux21_3 MUXNPC ( .a(NPCFromDecode), .b(OUT1RF), .sel(Mux1Sel), .y(MUXNPCout)
         );
  Mux21_2 MUXWITH4 ( .a({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b(MUX2out), .sel(Mux1Sel), .y(MUXWITH4out) );
  ALU_M32_C4 ALUset ( .CODE(ALUCODE), .DATA1(MUXNPCout), .DATA2(MUXWITH4out), 
        .OUTALU(ALUout) );
  reg_6 ALUout_REG ( .clock(clock), .reset(reset), .load(en3), .i(ALUout), .o(
        ALUtoMEMORY) );
  reg_5 RFout2_REG ( .clock(clock), .reset(reset), .load(en3), .i(OUT2RF), .o(
        OUT2RFtoMEMORY) );
  reg_4 AddressW_REG ( .clock(clock), .reset(reset), .load(en3), .i(
        AddressWfromDecode), .o(AddressWtoMEMORY) );
endmodule


module reg_3 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n215), .Z(n177) );
  BUF_X1 U4 ( .A(n215), .Z(n176) );
  BUF_X1 U5 ( .A(n215), .Z(n178) );
  BUF_X1 U6 ( .A(n216), .Z(n179) );
  BUF_X1 U7 ( .A(n216), .Z(n180) );
  BUF_X1 U8 ( .A(n216), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n215) );
  OAI22_X1 U10 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U12 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n213) );
  OAI22_X1 U14 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U16 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U18 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U20 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U22 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U24 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U26 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U28 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n205) );
  OAI22_X1 U30 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U32 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U34 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U36 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U38 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U40 ( .A1(n180), .A2(n51), .B1(n177), .B2(n199), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n199) );
  OAI22_X1 U42 ( .A1(n180), .A2(n52), .B1(n177), .B2(n198), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n198) );
  OAI22_X1 U44 ( .A1(n180), .A2(n53), .B1(n177), .B2(n197), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n197) );
  OAI22_X1 U46 ( .A1(n180), .A2(n54), .B1(n177), .B2(n196), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n196) );
  OAI22_X1 U48 ( .A1(n180), .A2(n55), .B1(n177), .B2(n195), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n195) );
  OAI22_X1 U50 ( .A1(n179), .A2(n56), .B1(n176), .B2(n194), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n194) );
  OAI22_X1 U52 ( .A1(n179), .A2(n57), .B1(n176), .B2(n193), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n193) );
  OAI22_X1 U54 ( .A1(n179), .A2(n58), .B1(n176), .B2(n192), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n192) );
  OAI22_X1 U56 ( .A1(n179), .A2(n59), .B1(n176), .B2(n191), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n191) );
  OAI22_X1 U58 ( .A1(n179), .A2(n60), .B1(n176), .B2(n190), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n190) );
  OAI22_X1 U60 ( .A1(n179), .A2(n61), .B1(n176), .B2(n189), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n189) );
  OAI22_X1 U62 ( .A1(n179), .A2(n62), .B1(n176), .B2(n188), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n188) );
  OAI22_X1 U64 ( .A1(n179), .A2(n63), .B1(n176), .B2(n187), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n187) );
  OAI22_X1 U66 ( .A1(n179), .A2(n64), .B1(n176), .B2(n186), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n186) );
  OAI22_X1 U68 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U70 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U72 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n183) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n216) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module reg_2 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n215), .Z(n177) );
  BUF_X1 U4 ( .A(n215), .Z(n176) );
  BUF_X1 U5 ( .A(n215), .Z(n178) );
  BUF_X1 U6 ( .A(n216), .Z(n179) );
  BUF_X1 U7 ( .A(n216), .Z(n180) );
  BUF_X1 U8 ( .A(n216), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n215) );
  OAI22_X1 U10 ( .A1(n181), .A2(n36), .B1(n178), .B2(n204), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n204) );
  OAI22_X1 U12 ( .A1(n181), .A2(n37), .B1(n178), .B2(n209), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n209) );
  OAI22_X1 U14 ( .A1(n181), .A2(n38), .B1(n178), .B2(n203), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n203) );
  OAI22_X1 U16 ( .A1(n181), .A2(n39), .B1(n178), .B2(n207), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n207) );
  OAI22_X1 U18 ( .A1(n181), .A2(n40), .B1(n178), .B2(n202), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n202) );
  OAI22_X1 U20 ( .A1(n181), .A2(n41), .B1(n178), .B2(n201), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n201) );
  OAI22_X1 U22 ( .A1(n181), .A2(n42), .B1(n178), .B2(n200), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n200) );
  OAI22_X1 U24 ( .A1(n180), .A2(n43), .B1(n178), .B2(n199), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n199) );
  OAI22_X1 U26 ( .A1(n180), .A2(n44), .B1(n177), .B2(n198), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n198) );
  OAI22_X1 U28 ( .A1(n180), .A2(n45), .B1(n177), .B2(n210), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n210) );
  OAI22_X1 U30 ( .A1(n180), .A2(n46), .B1(n177), .B2(n197), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n197) );
  OAI22_X1 U32 ( .A1(n180), .A2(n47), .B1(n177), .B2(n196), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n196) );
  OAI22_X1 U34 ( .A1(n180), .A2(n48), .B1(n177), .B2(n214), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n214) );
  OAI22_X1 U36 ( .A1(n180), .A2(n49), .B1(n177), .B2(n208), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n208) );
  OAI22_X1 U38 ( .A1(n180), .A2(n50), .B1(n177), .B2(n195), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n195) );
  OAI22_X1 U40 ( .A1(n180), .A2(n51), .B1(n177), .B2(n194), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n194) );
  OAI22_X1 U42 ( .A1(n180), .A2(n52), .B1(n177), .B2(n193), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n193) );
  OAI22_X1 U44 ( .A1(n180), .A2(n53), .B1(n177), .B2(n192), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n192) );
  OAI22_X1 U46 ( .A1(n180), .A2(n54), .B1(n177), .B2(n191), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n191) );
  OAI22_X1 U48 ( .A1(n180), .A2(n55), .B1(n177), .B2(n213), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n213) );
  OAI22_X1 U50 ( .A1(n179), .A2(n56), .B1(n176), .B2(n211), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n211) );
  OAI22_X1 U52 ( .A1(n179), .A2(n57), .B1(n176), .B2(n190), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n190) );
  OAI22_X1 U54 ( .A1(n179), .A2(n58), .B1(n176), .B2(n189), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n189) );
  OAI22_X1 U56 ( .A1(n179), .A2(n59), .B1(n176), .B2(n205), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n205) );
  OAI22_X1 U58 ( .A1(n179), .A2(n60), .B1(n176), .B2(n188), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n188) );
  OAI22_X1 U60 ( .A1(n179), .A2(n61), .B1(n176), .B2(n206), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n206) );
  OAI22_X1 U62 ( .A1(n179), .A2(n62), .B1(n176), .B2(n187), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n187) );
  OAI22_X1 U64 ( .A1(n179), .A2(n63), .B1(n176), .B2(n186), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n186) );
  OAI22_X1 U66 ( .A1(n179), .A2(n64), .B1(n176), .B2(n212), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n212) );
  OAI22_X1 U68 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U70 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U72 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n183) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n216) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module reg_1 ( clock, reset, load, i, o );
  input [31:0] i;
  output [31:0] o;
  input clock, reset, load;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216;

  DFF_X1 \temp_reg[31]  ( .D(n68), .CK(clock), .Q(o[31]), .QN(n67) );
  DFF_X1 \temp_reg[30]  ( .D(n69), .CK(clock), .Q(o[30]), .QN(n66) );
  DFF_X1 \temp_reg[29]  ( .D(n70), .CK(clock), .Q(o[29]), .QN(n65) );
  DFF_X1 \temp_reg[28]  ( .D(n71), .CK(clock), .Q(o[28]), .QN(n64) );
  DFF_X1 \temp_reg[27]  ( .D(n72), .CK(clock), .Q(o[27]), .QN(n63) );
  DFF_X1 \temp_reg[26]  ( .D(n73), .CK(clock), .Q(o[26]), .QN(n62) );
  DFF_X1 \temp_reg[25]  ( .D(n74), .CK(clock), .Q(o[25]), .QN(n61) );
  DFF_X1 \temp_reg[24]  ( .D(n75), .CK(clock), .Q(o[24]), .QN(n60) );
  DFF_X1 \temp_reg[23]  ( .D(n76), .CK(clock), .Q(o[23]), .QN(n59) );
  DFF_X1 \temp_reg[22]  ( .D(n77), .CK(clock), .Q(o[22]), .QN(n58) );
  DFF_X1 \temp_reg[21]  ( .D(n78), .CK(clock), .Q(o[21]), .QN(n57) );
  DFF_X1 \temp_reg[20]  ( .D(n79), .CK(clock), .Q(o[20]), .QN(n56) );
  DFF_X1 \temp_reg[19]  ( .D(n80), .CK(clock), .Q(o[19]), .QN(n55) );
  DFF_X1 \temp_reg[18]  ( .D(n81), .CK(clock), .Q(o[18]), .QN(n54) );
  DFF_X1 \temp_reg[17]  ( .D(n82), .CK(clock), .Q(o[17]), .QN(n53) );
  DFF_X1 \temp_reg[16]  ( .D(n83), .CK(clock), .Q(o[16]), .QN(n52) );
  DFF_X1 \temp_reg[15]  ( .D(n84), .CK(clock), .Q(o[15]), .QN(n51) );
  DFF_X1 \temp_reg[14]  ( .D(n85), .CK(clock), .Q(o[14]), .QN(n50) );
  DFF_X1 \temp_reg[13]  ( .D(n86), .CK(clock), .Q(o[13]), .QN(n49) );
  DFF_X1 \temp_reg[12]  ( .D(n87), .CK(clock), .Q(o[12]), .QN(n48) );
  DFF_X1 \temp_reg[11]  ( .D(n88), .CK(clock), .Q(o[11]), .QN(n47) );
  DFF_X1 \temp_reg[10]  ( .D(n89), .CK(clock), .Q(o[10]), .QN(n46) );
  DFF_X1 \temp_reg[9]  ( .D(n90), .CK(clock), .Q(o[9]), .QN(n45) );
  DFF_X1 \temp_reg[8]  ( .D(n91), .CK(clock), .Q(o[8]), .QN(n44) );
  DFF_X1 \temp_reg[7]  ( .D(n92), .CK(clock), .Q(o[7]), .QN(n43) );
  DFF_X1 \temp_reg[6]  ( .D(n93), .CK(clock), .Q(o[6]), .QN(n42) );
  DFF_X1 \temp_reg[5]  ( .D(n94), .CK(clock), .Q(o[5]), .QN(n41) );
  DFF_X1 \temp_reg[4]  ( .D(n95), .CK(clock), .Q(o[4]), .QN(n40) );
  DFF_X1 \temp_reg[3]  ( .D(n96), .CK(clock), .Q(o[3]), .QN(n39) );
  DFF_X1 \temp_reg[2]  ( .D(n97), .CK(clock), .Q(o[2]), .QN(n38) );
  DFF_X1 \temp_reg[1]  ( .D(n98), .CK(clock), .Q(o[1]), .QN(n37) );
  DFF_X1 \temp_reg[0]  ( .D(n99), .CK(clock), .Q(o[0]), .QN(n36) );
  BUF_X1 U3 ( .A(n215), .Z(n177) );
  BUF_X1 U4 ( .A(n215), .Z(n176) );
  BUF_X1 U5 ( .A(n215), .Z(n178) );
  BUF_X1 U6 ( .A(n216), .Z(n179) );
  BUF_X1 U7 ( .A(n216), .Z(n180) );
  BUF_X1 U8 ( .A(n216), .Z(n181) );
  NAND2_X1 U9 ( .A1(n182), .A2(n179), .ZN(n215) );
  OAI22_X1 U10 ( .A1(n181), .A2(n36), .B1(n178), .B2(n214), .ZN(n99) );
  INV_X1 U11 ( .A(i[0]), .ZN(n214) );
  OAI22_X1 U12 ( .A1(n181), .A2(n37), .B1(n178), .B2(n213), .ZN(n98) );
  INV_X1 U13 ( .A(i[1]), .ZN(n213) );
  OAI22_X1 U14 ( .A1(n181), .A2(n38), .B1(n178), .B2(n212), .ZN(n97) );
  INV_X1 U15 ( .A(i[2]), .ZN(n212) );
  OAI22_X1 U16 ( .A1(n181), .A2(n39), .B1(n178), .B2(n211), .ZN(n96) );
  INV_X1 U17 ( .A(i[3]), .ZN(n211) );
  OAI22_X1 U18 ( .A1(n181), .A2(n40), .B1(n178), .B2(n210), .ZN(n95) );
  INV_X1 U19 ( .A(i[4]), .ZN(n210) );
  OAI22_X1 U20 ( .A1(n181), .A2(n41), .B1(n178), .B2(n209), .ZN(n94) );
  INV_X1 U21 ( .A(i[5]), .ZN(n209) );
  OAI22_X1 U22 ( .A1(n181), .A2(n42), .B1(n178), .B2(n208), .ZN(n93) );
  INV_X1 U23 ( .A(i[6]), .ZN(n208) );
  OAI22_X1 U24 ( .A1(n180), .A2(n43), .B1(n178), .B2(n207), .ZN(n92) );
  INV_X1 U25 ( .A(i[7]), .ZN(n207) );
  OAI22_X1 U26 ( .A1(n180), .A2(n44), .B1(n177), .B2(n206), .ZN(n91) );
  INV_X1 U27 ( .A(i[8]), .ZN(n206) );
  OAI22_X1 U28 ( .A1(n180), .A2(n45), .B1(n177), .B2(n205), .ZN(n90) );
  INV_X1 U29 ( .A(i[9]), .ZN(n205) );
  OAI22_X1 U30 ( .A1(n180), .A2(n46), .B1(n177), .B2(n204), .ZN(n89) );
  INV_X1 U31 ( .A(i[10]), .ZN(n204) );
  OAI22_X1 U32 ( .A1(n180), .A2(n47), .B1(n177), .B2(n203), .ZN(n88) );
  INV_X1 U33 ( .A(i[11]), .ZN(n203) );
  OAI22_X1 U34 ( .A1(n180), .A2(n48), .B1(n177), .B2(n202), .ZN(n87) );
  INV_X1 U35 ( .A(i[12]), .ZN(n202) );
  OAI22_X1 U36 ( .A1(n180), .A2(n49), .B1(n177), .B2(n201), .ZN(n86) );
  INV_X1 U37 ( .A(i[13]), .ZN(n201) );
  OAI22_X1 U38 ( .A1(n180), .A2(n50), .B1(n177), .B2(n200), .ZN(n85) );
  INV_X1 U39 ( .A(i[14]), .ZN(n200) );
  OAI22_X1 U40 ( .A1(n180), .A2(n51), .B1(n177), .B2(n199), .ZN(n84) );
  INV_X1 U41 ( .A(i[15]), .ZN(n199) );
  OAI22_X1 U42 ( .A1(n180), .A2(n52), .B1(n177), .B2(n198), .ZN(n83) );
  INV_X1 U43 ( .A(i[16]), .ZN(n198) );
  OAI22_X1 U44 ( .A1(n180), .A2(n53), .B1(n177), .B2(n197), .ZN(n82) );
  INV_X1 U45 ( .A(i[17]), .ZN(n197) );
  OAI22_X1 U46 ( .A1(n180), .A2(n54), .B1(n177), .B2(n196), .ZN(n81) );
  INV_X1 U47 ( .A(i[18]), .ZN(n196) );
  OAI22_X1 U48 ( .A1(n180), .A2(n55), .B1(n177), .B2(n195), .ZN(n80) );
  INV_X1 U49 ( .A(i[19]), .ZN(n195) );
  OAI22_X1 U50 ( .A1(n179), .A2(n56), .B1(n176), .B2(n194), .ZN(n79) );
  INV_X1 U51 ( .A(i[20]), .ZN(n194) );
  OAI22_X1 U52 ( .A1(n179), .A2(n57), .B1(n176), .B2(n193), .ZN(n78) );
  INV_X1 U53 ( .A(i[21]), .ZN(n193) );
  OAI22_X1 U54 ( .A1(n179), .A2(n58), .B1(n176), .B2(n192), .ZN(n77) );
  INV_X1 U55 ( .A(i[22]), .ZN(n192) );
  OAI22_X1 U56 ( .A1(n179), .A2(n59), .B1(n176), .B2(n191), .ZN(n76) );
  INV_X1 U57 ( .A(i[23]), .ZN(n191) );
  OAI22_X1 U58 ( .A1(n179), .A2(n60), .B1(n176), .B2(n190), .ZN(n75) );
  INV_X1 U59 ( .A(i[24]), .ZN(n190) );
  OAI22_X1 U60 ( .A1(n179), .A2(n61), .B1(n176), .B2(n189), .ZN(n74) );
  INV_X1 U61 ( .A(i[25]), .ZN(n189) );
  OAI22_X1 U62 ( .A1(n179), .A2(n62), .B1(n176), .B2(n188), .ZN(n73) );
  INV_X1 U63 ( .A(i[26]), .ZN(n188) );
  OAI22_X1 U64 ( .A1(n179), .A2(n63), .B1(n176), .B2(n187), .ZN(n72) );
  INV_X1 U65 ( .A(i[27]), .ZN(n187) );
  OAI22_X1 U66 ( .A1(n179), .A2(n64), .B1(n176), .B2(n186), .ZN(n71) );
  INV_X1 U67 ( .A(i[28]), .ZN(n186) );
  OAI22_X1 U68 ( .A1(n179), .A2(n65), .B1(n176), .B2(n185), .ZN(n70) );
  INV_X1 U69 ( .A(i[29]), .ZN(n185) );
  OAI22_X1 U70 ( .A1(n179), .A2(n66), .B1(n176), .B2(n184), .ZN(n69) );
  INV_X1 U71 ( .A(i[30]), .ZN(n184) );
  OAI22_X1 U72 ( .A1(n179), .A2(n67), .B1(n176), .B2(n183), .ZN(n68) );
  INV_X1 U73 ( .A(i[31]), .ZN(n183) );
  OR2_X1 U74 ( .A1(load), .A2(reset), .ZN(n216) );
  INV_X1 U75 ( .A(reset), .ZN(n182) );
endmodule


module memoryUnit ( clock, reset, en4, ALUout, DRAMout, AddressWfromEXECUTE, 
        LOADDATA, ALUtoWBMUX, AddressWtoWB );
  input [31:0] ALUout;
  input [31:0] DRAMout;
  input [31:0] AddressWfromEXECUTE;
  output [31:0] LOADDATA;
  output [31:0] ALUtoWBMUX;
  output [31:0] AddressWtoWB;
  input clock, reset, en4;


  reg_3 LMD_REG ( .clock(clock), .reset(reset), .load(en4), .i(DRAMout), .o(
        LOADDATA) );
  reg_2 ALUout_REG ( .clock(clock), .reset(reset), .load(en4), .i(ALUout), .o(
        ALUtoWBMUX) );
  reg_1 AddressW_REG ( .clock(clock), .reset(reset), .load(en4), .i(
        AddressWfromEXECUTE), .o(AddressWtoWB) );
endmodule


module Mux21_1 ( a, b, sel, y );
  input [31:0] a;
  input [31:0] b;
  output [31:0] y;
  input sel;
  wire   n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246;

  INV_X1 U1 ( .A(n181), .ZN(n172) );
  BUF_X1 U2 ( .A(n182), .Z(n173) );
  BUF_X1 U3 ( .A(n173), .Z(n180) );
  BUF_X1 U4 ( .A(n175), .Z(n179) );
  BUF_X1 U5 ( .A(n182), .Z(n178) );
  BUF_X1 U6 ( .A(n182), .Z(n177) );
  BUF_X1 U7 ( .A(n182), .Z(n176) );
  BUF_X1 U8 ( .A(n182), .Z(n175) );
  BUF_X1 U9 ( .A(n182), .Z(n174) );
  BUF_X1 U10 ( .A(n182), .Z(n181) );
  INV_X1 U11 ( .A(sel), .ZN(n182) );
  INV_X1 U12 ( .A(n240), .ZN(y[3]) );
  AOI22_X1 U13 ( .A1(a[3]), .A2(n172), .B1(b[3]), .B2(n174), .ZN(n240) );
  INV_X1 U14 ( .A(n241), .ZN(y[4]) );
  AOI22_X1 U15 ( .A1(a[4]), .A2(n172), .B1(b[4]), .B2(n174), .ZN(n241) );
  INV_X1 U16 ( .A(n242), .ZN(y[5]) );
  AOI22_X1 U17 ( .A1(a[5]), .A2(n172), .B1(b[5]), .B2(n174), .ZN(n242) );
  INV_X1 U18 ( .A(n243), .ZN(y[6]) );
  AOI22_X1 U19 ( .A1(a[6]), .A2(n172), .B1(b[6]), .B2(n173), .ZN(n243) );
  INV_X1 U20 ( .A(n244), .ZN(y[7]) );
  AOI22_X1 U21 ( .A1(a[7]), .A2(n172), .B1(b[7]), .B2(n173), .ZN(n244) );
  INV_X1 U22 ( .A(n245), .ZN(y[8]) );
  AOI22_X1 U23 ( .A1(a[8]), .A2(n172), .B1(b[8]), .B2(n173), .ZN(n245) );
  INV_X1 U24 ( .A(n239), .ZN(y[31]) );
  AOI22_X1 U25 ( .A1(a[31]), .A2(sel), .B1(b[31]), .B2(n174), .ZN(n239) );
  INV_X1 U26 ( .A(n215), .ZN(y[0]) );
  AOI22_X1 U27 ( .A1(a[0]), .A2(n172), .B1(b[0]), .B2(n180), .ZN(n215) );
  INV_X1 U28 ( .A(n226), .ZN(y[1]) );
  AOI22_X1 U29 ( .A1(a[1]), .A2(n172), .B1(b[1]), .B2(n178), .ZN(n226) );
  INV_X1 U30 ( .A(n237), .ZN(y[2]) );
  AOI22_X1 U31 ( .A1(a[2]), .A2(sel), .B1(b[2]), .B2(n175), .ZN(n237) );
  INV_X1 U32 ( .A(n216), .ZN(y[10]) );
  AOI22_X1 U33 ( .A1(a[10]), .A2(n172), .B1(b[10]), .B2(n180), .ZN(n216) );
  INV_X1 U34 ( .A(n217), .ZN(y[11]) );
  AOI22_X1 U35 ( .A1(a[11]), .A2(n172), .B1(b[11]), .B2(n180), .ZN(n217) );
  INV_X1 U36 ( .A(n218), .ZN(y[12]) );
  AOI22_X1 U37 ( .A1(a[12]), .A2(n172), .B1(b[12]), .B2(n180), .ZN(n218) );
  INV_X1 U38 ( .A(n219), .ZN(y[13]) );
  AOI22_X1 U39 ( .A1(a[13]), .A2(n172), .B1(b[13]), .B2(n179), .ZN(n219) );
  INV_X1 U40 ( .A(n220), .ZN(y[14]) );
  AOI22_X1 U41 ( .A1(a[14]), .A2(n172), .B1(b[14]), .B2(n179), .ZN(n220) );
  INV_X1 U42 ( .A(n221), .ZN(y[15]) );
  AOI22_X1 U43 ( .A1(a[15]), .A2(n172), .B1(b[15]), .B2(n179), .ZN(n221) );
  INV_X1 U44 ( .A(n222), .ZN(y[16]) );
  AOI22_X1 U45 ( .A1(a[16]), .A2(n172), .B1(b[16]), .B2(n179), .ZN(n222) );
  INV_X1 U46 ( .A(n223), .ZN(y[17]) );
  AOI22_X1 U47 ( .A1(a[17]), .A2(n172), .B1(b[17]), .B2(n178), .ZN(n223) );
  INV_X1 U48 ( .A(n224), .ZN(y[18]) );
  AOI22_X1 U49 ( .A1(a[18]), .A2(n172), .B1(b[18]), .B2(n178), .ZN(n224) );
  INV_X1 U50 ( .A(n225), .ZN(y[19]) );
  AOI22_X1 U51 ( .A1(a[19]), .A2(n172), .B1(b[19]), .B2(n178), .ZN(n225) );
  INV_X1 U52 ( .A(n227), .ZN(y[20]) );
  AOI22_X1 U53 ( .A1(a[20]), .A2(sel), .B1(b[20]), .B2(n177), .ZN(n227) );
  INV_X1 U54 ( .A(n228), .ZN(y[21]) );
  AOI22_X1 U55 ( .A1(a[21]), .A2(sel), .B1(b[21]), .B2(n177), .ZN(n228) );
  INV_X1 U56 ( .A(n229), .ZN(y[22]) );
  AOI22_X1 U57 ( .A1(a[22]), .A2(sel), .B1(b[22]), .B2(n177), .ZN(n229) );
  INV_X1 U58 ( .A(n230), .ZN(y[23]) );
  AOI22_X1 U59 ( .A1(a[23]), .A2(sel), .B1(b[23]), .B2(n177), .ZN(n230) );
  INV_X1 U60 ( .A(n231), .ZN(y[24]) );
  AOI22_X1 U61 ( .A1(a[24]), .A2(sel), .B1(b[24]), .B2(n176), .ZN(n231) );
  INV_X1 U62 ( .A(n232), .ZN(y[25]) );
  AOI22_X1 U63 ( .A1(a[25]), .A2(sel), .B1(b[25]), .B2(n176), .ZN(n232) );
  INV_X1 U64 ( .A(n233), .ZN(y[26]) );
  AOI22_X1 U65 ( .A1(a[26]), .A2(sel), .B1(b[26]), .B2(n176), .ZN(n233) );
  INV_X1 U66 ( .A(n234), .ZN(y[27]) );
  AOI22_X1 U67 ( .A1(a[27]), .A2(sel), .B1(b[27]), .B2(n176), .ZN(n234) );
  INV_X1 U68 ( .A(n235), .ZN(y[28]) );
  AOI22_X1 U69 ( .A1(a[28]), .A2(sel), .B1(b[28]), .B2(n175), .ZN(n235) );
  INV_X1 U70 ( .A(n236), .ZN(y[29]) );
  AOI22_X1 U71 ( .A1(a[29]), .A2(sel), .B1(b[29]), .B2(n175), .ZN(n236) );
  INV_X1 U72 ( .A(n238), .ZN(y[30]) );
  AOI22_X1 U73 ( .A1(a[30]), .A2(sel), .B1(b[30]), .B2(n175), .ZN(n238) );
  INV_X1 U74 ( .A(n246), .ZN(y[9]) );
  AOI22_X1 U75 ( .A1(sel), .A2(a[9]), .B1(b[9]), .B2(n173), .ZN(n246) );
endmodule


module WBUnit ( selwb, ALUin, LOADDATA, AddressWfromMemory, MUXtoRF, 
        AddressWtoDECODE );
  input [31:0] ALUin;
  input [31:0] LOADDATA;
  input [31:0] AddressWfromMemory;
  output [31:0] MUXtoRF;
  output [31:0] AddressWtoDECODE;
  input selwb;

  assign AddressWtoDECODE[31] = AddressWfromMemory[31];
  assign AddressWtoDECODE[30] = AddressWfromMemory[30];
  assign AddressWtoDECODE[29] = AddressWfromMemory[29];
  assign AddressWtoDECODE[28] = AddressWfromMemory[28];
  assign AddressWtoDECODE[27] = AddressWfromMemory[27];
  assign AddressWtoDECODE[26] = AddressWfromMemory[26];
  assign AddressWtoDECODE[25] = AddressWfromMemory[25];
  assign AddressWtoDECODE[24] = AddressWfromMemory[24];
  assign AddressWtoDECODE[23] = AddressWfromMemory[23];
  assign AddressWtoDECODE[22] = AddressWfromMemory[22];
  assign AddressWtoDECODE[21] = AddressWfromMemory[21];
  assign AddressWtoDECODE[20] = AddressWfromMemory[20];
  assign AddressWtoDECODE[19] = AddressWfromMemory[19];
  assign AddressWtoDECODE[18] = AddressWfromMemory[18];
  assign AddressWtoDECODE[17] = AddressWfromMemory[17];
  assign AddressWtoDECODE[16] = AddressWfromMemory[16];
  assign AddressWtoDECODE[15] = AddressWfromMemory[15];
  assign AddressWtoDECODE[14] = AddressWfromMemory[14];
  assign AddressWtoDECODE[13] = AddressWfromMemory[13];
  assign AddressWtoDECODE[12] = AddressWfromMemory[12];
  assign AddressWtoDECODE[11] = AddressWfromMemory[11];
  assign AddressWtoDECODE[10] = AddressWfromMemory[10];
  assign AddressWtoDECODE[9] = AddressWfromMemory[9];
  assign AddressWtoDECODE[8] = AddressWfromMemory[8];
  assign AddressWtoDECODE[7] = AddressWfromMemory[7];
  assign AddressWtoDECODE[6] = AddressWfromMemory[6];
  assign AddressWtoDECODE[5] = AddressWfromMemory[5];
  assign AddressWtoDECODE[4] = AddressWfromMemory[4];
  assign AddressWtoDECODE[3] = AddressWfromMemory[3];
  assign AddressWtoDECODE[2] = AddressWfromMemory[2];
  assign AddressWtoDECODE[1] = AddressWfromMemory[1];
  assign AddressWtoDECODE[0] = AddressWfromMemory[0];

  Mux21_1 wbmux ( .a(LOADDATA), .b(ALUin), .sel(selwb), .y(MUXtoRF) );
endmodule


module dataPath_M32_C4_N5 ( clock, reset, Instruction, en1, en2, SignSelect, 
        RD1, RD2, WR, JMP, BRANCHenable, en3, BranchCondSel, Mux1Sel, Mux2Sel, 
        ALUCODE, RegDestination, en4, DRAMout, selwb, PCtoIM, ALUtoMEMORY, 
        OUT2RFtoMEMORY, InstructionToCU );
  input [31:0] Instruction;
  input [3:0] ALUCODE;
  input [31:0] DRAMout;
  output [31:0] PCtoIM;
  output [31:0] ALUtoMEMORY;
  output [31:0] OUT2RFtoMEMORY;
  output [31:0] InstructionToCU;
  input clock, reset, en1, en2, SignSelect, RD1, RD2, WR, JMP, BRANCHenable,
         en3, BranchCondSel, Mux1Sel, Mux2Sel, RegDestination, en4, selwb;
  wire   BRANCHtoFetch, n1;
  wire   [31:0] NewPC;
  wire   [31:0] NXPC;
  wire   [4:0] AddressfromWB;
  wire   [31:0] MUXtoRF;
  wire   [31:0] OUT1;
  wire   [31:0] OUT2;
  wire   [31:0] OUTIMM;
  wire   [31:0] NPCfromDECODE;
  wire   [31:0] ADDWfromDECODE;
  wire   [31:0] ADDWtoMEMORY;
  wire   [31:0] LOADDATA;
  wire   [31:0] ALUtoWBMUX;
  wire   [31:0] ADDWtoWB;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48;

  fetchUnit FU ( .clock(clock), .reset(n1), .en1(en1), .BranchPC({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, NewPC[9:0]}), 
        .BRANCHfromDECODE(BRANCHtoFetch), .Instruction(Instruction), .PCtoIM(
        PCtoIM), .IRtoDecode(InstructionToCU), .NPCtoDecode(NXPC) );
  DecodeUnit DU ( .clock(clock), .reset(n1), .JMP(JMP), .RegDestination(
        RegDestination), .en2(en2), .SignSelect(SignSelect), .BranchCondSel(
        BranchCondSel), .BRANCHenable(BRANCHenable), .RD1(RD1), .RD2(RD2), 
        .WR(WR), .Instruction(InstructionToCU), .ADD_WR(AddressfromWB), 
        .DATAIN(MUXtoRF), .NPCfromIF(NXPC), .OUT1(OUT1), .OUT2(OUT2), .OUTNPC(
        {SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, NewPC[9:0]}), 
        .OUTIMM(OUTIMM), .NPCtoEX(NPCfromDECODE), .AddressWtoEX(ADDWfromDECODE), .BRANCHtoFetch(BRANCHtoFetch) );
  executeUnit_M32_C4 EU ( .clock(clock), .reset(n1), .en3(en3), .Mux1Sel(
        Mux1Sel), .Mux2Sel(Mux2Sel), .ALUCODE(ALUCODE), .OUT1RF(OUT1), 
        .OUT2RF(OUT2), .IMMEDIATE(OUTIMM), .NPCFromDecode(NPCfromDECODE), 
        .AddressWfromDecode(ADDWfromDECODE), .ALUtoMEMORY(ALUtoMEMORY), 
        .OUT2RFtoMEMORY(OUT2RFtoMEMORY), .AddressWtoMEMORY(ADDWtoMEMORY) );
  memoryUnit MU ( .clock(clock), .reset(n1), .en4(en4), .ALUout(ALUtoMEMORY), 
        .DRAMout(DRAMout), .AddressWfromEXECUTE(ADDWtoMEMORY), .LOADDATA(
        LOADDATA), .ALUtoWBMUX(ALUtoWBMUX), .AddressWtoWB(ADDWtoWB) );
  WBUnit WBU ( .selwb(selwb), .ALUin(ALUtoWBMUX), .LOADDATA(LOADDATA), 
        .AddressWfromMemory(ADDWtoWB), .MUXtoRF(MUXtoRF), .AddressWtoDECODE({
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, AddressfromWB}) );
  BUF_X1 U23 ( .A(reset), .Z(n1) );
endmodule


module DLX_M32_C4_N5 ( Clk, Rst, IRAM_Addr, IRAM_Dout, DRAM_MemoryEnable, 
        DRAM_ReadNotWrite, DRAM_Addr, DRAM_in, DRAM_out );
  output [31:0] IRAM_Addr;
  input [31:0] IRAM_Dout;
  output [4:0] DRAM_Addr;
  output [31:0] DRAM_in;
  input [31:0] DRAM_out;
  input Clk, Rst;
  output DRAM_MemoryEnable, DRAM_ReadNotWrite;
  wire   en2, SignSelect, RD1, RD2, JMP, BranchCondSel, BRANCHenable,
         RegDestination, en3, Mux1Sel, Mux2Sel, en4, selwb, WR;
  wire   [31:0] InstructionToCU;
  wire   [3:0] ALUCODE;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26;

  Cu_M32_FUNC_SIZE11_OP_CODE_SIZE6_ALU_OP_CODE_SIZE4_CW_SIZE17 CU_I ( .Clk(Clk), .Rst(Rst), .IR_IN(InstructionToCU), .en2(en2), .SignSelect(SignSelect), 
        .RD1(RD1), .RD2(RD2), .JMP(JMP), .BranchCondSel(BranchCondSel), 
        .BRANCHenable(BRANCHenable), .RegDestination(RegDestination), .en3(en3), .Mux1Sel(Mux1Sel), .Mux2Sel(Mux2Sel), .ALUCODE(ALUCODE), .en4(en4), 
        .MemoryEnable(DRAM_MemoryEnable), .ReadNotWrite(DRAM_ReadNotWrite), 
        .selwb(selwb), .WR(WR) );
  dataPath_M32_C4_N5 DP ( .clock(Clk), .reset(Rst), .Instruction(IRAM_Dout), 
        .en1(1'b1), .en2(en2), .SignSelect(SignSelect), .RD1(RD1), .RD2(RD2), 
        .WR(WR), .JMP(JMP), .BRANCHenable(BRANCHenable), .en3(en3), 
        .BranchCondSel(BranchCondSel), .Mux1Sel(Mux1Sel), .Mux2Sel(Mux2Sel), 
        .ALUCODE(ALUCODE), .RegDestination(RegDestination), .en4(en4), 
        .DRAMout(DRAM_out), .selwb(selwb), .PCtoIM(IRAM_Addr), .ALUtoMEMORY({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, DRAM_Addr}), .OUT2RFtoMEMORY(DRAM_in), 
        .InstructionToCU(InstructionToCU) );
endmodule

